module lpif_txrx_x16_h2_master_concat  (

// Data from Logic Links
  input  logic [ 588:   0]   tx_downstream_data  ,
  output logic               tx_downstream_pop_ovrd,

  output logic [ 588:   0]   rx_upstream_data    ,
  output logic               rx_upstream_push_ovrd,

// PHY Interconnect
  output logic [ 159:   0]   tx_phy0             ,
  input  logic [ 159:   0]   rx_phy0             ,
  output logic [ 159:   0]   tx_phy1             ,
  input  logic [ 159:   0]   rx_phy1             ,
  output logic [ 159:   0]   tx_phy2             ,
  input  logic [ 159:   0]   rx_phy2             ,
  output logic [ 159:   0]   tx_phy3             ,
  input  logic [ 159:   0]   rx_phy3             ,

  input  logic               clk_wr              ,
  input  logic               clk_rd              ,
  input  logic               rst_wr_n            ,
  input  logic               rst_rd_n            ,

  input  logic               m_gen2_mode         ,
  input  logic               tx_online           ,

  input  logic               tx_stb_userbit      ,
  input  logic [   1:   0]   tx_mrk_userbit      

);

// No TX Packetization, so tie off packetization signals
  assign tx_downstream_pop_ovrd               = 1'b0                               ;

// No RX Packetization, so tie off packetization signals
  assign rx_upstream_push_ovrd               = 1'b0                               ;

//////////////////////////////////////////////////////////////////
// TX Section

//   TX_CH_WIDTH           = 160; // Gen2 running at Half Rate
//   TX_DATA_WIDTH         = 157; // Usable Data per Channel
//   TX_PERSISTENT_STROBE  = 1'b1;
//   TX_PERSISTENT_MARKER  = 1'b1;
//   TX_STROBE_GEN2_LOC    = 'd76;
//   TX_MARKER_GEN2_LOC    = 'd4;
//   TX_STROBE_GEN1_LOC    = 'd38;
//   TX_MARKER_GEN1_LOC    = 'd39;
//   TX_ENABLE_STROBE      = 1'b1;
//   TX_ENABLE_MARKER      = 1'b1;
//   TX_DBI_PRESENT        = 1'b0;
//   TX_REG_PHY            = 1'b0;

  localparam TX_REG_PHY    = 1'b0;  // If set, this enables boundary FF for timing reasons

  logic [ 159:   0]                              tx_phy_preflop_0              ;
  logic [ 159:   0]                              tx_phy_preflop_1              ;
  logic [ 159:   0]                              tx_phy_preflop_2              ;
  logic [ 159:   0]                              tx_phy_preflop_3              ;
  logic [ 159:   0]                              tx_phy_flop_0_reg             ;
  logic [ 159:   0]                              tx_phy_flop_1_reg             ;
  logic [ 159:   0]                              tx_phy_flop_2_reg             ;
  logic [ 159:   0]                              tx_phy_flop_3_reg             ;

  always_ff @(posedge clk_wr or negedge rst_wr_n)
  if (~rst_wr_n)
  begin
    tx_phy_flop_0_reg                       <= 160'b0                                  ;
    tx_phy_flop_1_reg                       <= 160'b0                                  ;
    tx_phy_flop_2_reg                       <= 160'b0                                  ;
    tx_phy_flop_3_reg                       <= 160'b0                                  ;
  end
  else
  begin
    tx_phy_flop_0_reg                       <= tx_phy_preflop_0                        ;
    tx_phy_flop_1_reg                       <= tx_phy_preflop_1                        ;
    tx_phy_flop_2_reg                       <= tx_phy_preflop_2                        ;
    tx_phy_flop_3_reg                       <= tx_phy_preflop_3                        ;
  end

  assign tx_phy0                            = TX_REG_PHY ? tx_phy_flop_0_reg : tx_phy_preflop_0               ;
  assign tx_phy1                            = TX_REG_PHY ? tx_phy_flop_1_reg : tx_phy_preflop_1               ;
  assign tx_phy2                            = TX_REG_PHY ? tx_phy_flop_2_reg : tx_phy_preflop_2               ;
  assign tx_phy3                            = TX_REG_PHY ? tx_phy_flop_3_reg : tx_phy_preflop_3               ;

  assign tx_phy_preflop_0 [   0] = tx_downstream_data  [   0] ;
  assign tx_phy_preflop_0 [   1] = tx_downstream_data  [   1] ;
  assign tx_phy_preflop_0 [   2] = tx_downstream_data  [   2] ;
  assign tx_phy_preflop_0 [   3] = tx_downstream_data  [   3] ;
  assign tx_phy_preflop_0 [   4] = tx_mrk_userbit[0]          ; // MARKER
  assign tx_phy_preflop_0 [   5] = tx_downstream_data  [   4] ;
  assign tx_phy_preflop_0 [   6] = tx_downstream_data  [   5] ;
  assign tx_phy_preflop_0 [   7] = tx_downstream_data  [   6] ;
  assign tx_phy_preflop_0 [   8] = tx_downstream_data  [   7] ;
  assign tx_phy_preflop_0 [   9] = tx_downstream_data  [   8] ;
  assign tx_phy_preflop_0 [  10] = tx_downstream_data  [   9] ;
  assign tx_phy_preflop_0 [  11] = tx_downstream_data  [  10] ;
  assign tx_phy_preflop_0 [  12] = tx_downstream_data  [  11] ;
  assign tx_phy_preflop_0 [  13] = tx_downstream_data  [  12] ;
  assign tx_phy_preflop_0 [  14] = tx_downstream_data  [  13] ;
  assign tx_phy_preflop_0 [  15] = tx_downstream_data  [  14] ;
  assign tx_phy_preflop_0 [  16] = tx_downstream_data  [  15] ;
  assign tx_phy_preflop_0 [  17] = tx_downstream_data  [  16] ;
  assign tx_phy_preflop_0 [  18] = tx_downstream_data  [  17] ;
  assign tx_phy_preflop_0 [  19] = tx_downstream_data  [  18] ;
  assign tx_phy_preflop_0 [  20] = tx_downstream_data  [  19] ;
  assign tx_phy_preflop_0 [  21] = tx_downstream_data  [  20] ;
  assign tx_phy_preflop_0 [  22] = tx_downstream_data  [  21] ;
  assign tx_phy_preflop_0 [  23] = tx_downstream_data  [  22] ;
  assign tx_phy_preflop_0 [  24] = tx_downstream_data  [  23] ;
  assign tx_phy_preflop_0 [  25] = tx_downstream_data  [  24] ;
  assign tx_phy_preflop_0 [  26] = tx_downstream_data  [  25] ;
  assign tx_phy_preflop_0 [  27] = tx_downstream_data  [  26] ;
  assign tx_phy_preflop_0 [  28] = tx_downstream_data  [  27] ;
  assign tx_phy_preflop_0 [  29] = tx_downstream_data  [  28] ;
  assign tx_phy_preflop_0 [  30] = tx_downstream_data  [  29] ;
  assign tx_phy_preflop_0 [  31] = tx_downstream_data  [  30] ;
  assign tx_phy_preflop_0 [  32] = tx_downstream_data  [  31] ;
  assign tx_phy_preflop_0 [  33] = tx_downstream_data  [  32] ;
  assign tx_phy_preflop_0 [  34] = tx_downstream_data  [  33] ;
  assign tx_phy_preflop_0 [  35] = tx_downstream_data  [  34] ;
  assign tx_phy_preflop_0 [  36] = tx_downstream_data  [  35] ;
  assign tx_phy_preflop_0 [  37] = tx_downstream_data  [  36] ;
  assign tx_phy_preflop_0 [  38] = tx_downstream_data  [  37] ;
  assign tx_phy_preflop_0 [  39] = tx_downstream_data  [  38] ;
  assign tx_phy_preflop_0 [  40] = tx_downstream_data  [  39] ;
  assign tx_phy_preflop_0 [  41] = tx_downstream_data  [  40] ;
  assign tx_phy_preflop_0 [  42] = tx_downstream_data  [  41] ;
  assign tx_phy_preflop_0 [  43] = tx_downstream_data  [  42] ;
  assign tx_phy_preflop_0 [  44] = tx_downstream_data  [  43] ;
  assign tx_phy_preflop_0 [  45] = tx_downstream_data  [  44] ;
  assign tx_phy_preflop_0 [  46] = tx_downstream_data  [  45] ;
  assign tx_phy_preflop_0 [  47] = tx_downstream_data  [  46] ;
  assign tx_phy_preflop_0 [  48] = tx_downstream_data  [  47] ;
  assign tx_phy_preflop_0 [  49] = tx_downstream_data  [  48] ;
  assign tx_phy_preflop_0 [  50] = tx_downstream_data  [  49] ;
  assign tx_phy_preflop_0 [  51] = tx_downstream_data  [  50] ;
  assign tx_phy_preflop_0 [  52] = tx_downstream_data  [  51] ;
  assign tx_phy_preflop_0 [  53] = tx_downstream_data  [  52] ;
  assign tx_phy_preflop_0 [  54] = tx_downstream_data  [  53] ;
  assign tx_phy_preflop_0 [  55] = tx_downstream_data  [  54] ;
  assign tx_phy_preflop_0 [  56] = tx_downstream_data  [  55] ;
  assign tx_phy_preflop_0 [  57] = tx_downstream_data  [  56] ;
  assign tx_phy_preflop_0 [  58] = tx_downstream_data  [  57] ;
  assign tx_phy_preflop_0 [  59] = tx_downstream_data  [  58] ;
  assign tx_phy_preflop_0 [  60] = tx_downstream_data  [  59] ;
  assign tx_phy_preflop_0 [  61] = tx_downstream_data  [  60] ;
  assign tx_phy_preflop_0 [  62] = tx_downstream_data  [  61] ;
  assign tx_phy_preflop_0 [  63] = tx_downstream_data  [  62] ;
  assign tx_phy_preflop_0 [  64] = tx_downstream_data  [  63] ;
  assign tx_phy_preflop_0 [  65] = tx_downstream_data  [  64] ;
  assign tx_phy_preflop_0 [  66] = tx_downstream_data  [  65] ;
  assign tx_phy_preflop_0 [  67] = tx_downstream_data  [  66] ;
  assign tx_phy_preflop_0 [  68] = tx_downstream_data  [  67] ;
  assign tx_phy_preflop_0 [  69] = tx_downstream_data  [  68] ;
  assign tx_phy_preflop_0 [  70] = tx_downstream_data  [  69] ;
  assign tx_phy_preflop_0 [  71] = tx_downstream_data  [  70] ;
  assign tx_phy_preflop_0 [  72] = tx_downstream_data  [  71] ;
  assign tx_phy_preflop_0 [  73] = tx_downstream_data  [  72] ;
  assign tx_phy_preflop_0 [  74] = tx_downstream_data  [  73] ;
  assign tx_phy_preflop_0 [  75] = tx_downstream_data  [  74] ;
  assign tx_phy_preflop_0 [  76] = tx_stb_userbit             ; // STROBE
  assign tx_phy_preflop_0 [  77] = tx_downstream_data  [  75] ;
  assign tx_phy_preflop_0 [  78] = tx_downstream_data  [  76] ;
  assign tx_phy_preflop_0 [  79] = tx_downstream_data  [  77] ;
  assign tx_phy_preflop_0 [  80] = tx_downstream_data  [  78] ;
  assign tx_phy_preflop_0 [  81] = tx_downstream_data  [  79] ;
  assign tx_phy_preflop_0 [  82] = tx_downstream_data  [  80] ;
  assign tx_phy_preflop_0 [  83] = tx_downstream_data  [  81] ;
  assign tx_phy_preflop_0 [  84] = tx_mrk_userbit[1]          ; // MARKER
  assign tx_phy_preflop_0 [  85] = tx_downstream_data  [  82] ;
  assign tx_phy_preflop_0 [  86] = tx_downstream_data  [  83] ;
  assign tx_phy_preflop_0 [  87] = tx_downstream_data  [  84] ;
  assign tx_phy_preflop_0 [  88] = tx_downstream_data  [  85] ;
  assign tx_phy_preflop_0 [  89] = tx_downstream_data  [  86] ;
  assign tx_phy_preflop_0 [  90] = tx_downstream_data  [  87] ;
  assign tx_phy_preflop_0 [  91] = tx_downstream_data  [  88] ;
  assign tx_phy_preflop_0 [  92] = tx_downstream_data  [  89] ;
  assign tx_phy_preflop_0 [  93] = tx_downstream_data  [  90] ;
  assign tx_phy_preflop_0 [  94] = tx_downstream_data  [  91] ;
  assign tx_phy_preflop_0 [  95] = tx_downstream_data  [  92] ;
  assign tx_phy_preflop_0 [  96] = tx_downstream_data  [  93] ;
  assign tx_phy_preflop_0 [  97] = tx_downstream_data  [  94] ;
  assign tx_phy_preflop_0 [  98] = tx_downstream_data  [  95] ;
  assign tx_phy_preflop_0 [  99] = tx_downstream_data  [  96] ;
  assign tx_phy_preflop_0 [ 100] = tx_downstream_data  [  97] ;
  assign tx_phy_preflop_0 [ 101] = tx_downstream_data  [  98] ;
  assign tx_phy_preflop_0 [ 102] = tx_downstream_data  [  99] ;
  assign tx_phy_preflop_0 [ 103] = tx_downstream_data  [ 100] ;
  assign tx_phy_preflop_0 [ 104] = tx_downstream_data  [ 101] ;
  assign tx_phy_preflop_0 [ 105] = tx_downstream_data  [ 102] ;
  assign tx_phy_preflop_0 [ 106] = tx_downstream_data  [ 103] ;
  assign tx_phy_preflop_0 [ 107] = tx_downstream_data  [ 104] ;
  assign tx_phy_preflop_0 [ 108] = tx_downstream_data  [ 105] ;
  assign tx_phy_preflop_0 [ 109] = tx_downstream_data  [ 106] ;
  assign tx_phy_preflop_0 [ 110] = tx_downstream_data  [ 107] ;
  assign tx_phy_preflop_0 [ 111] = tx_downstream_data  [ 108] ;
  assign tx_phy_preflop_0 [ 112] = tx_downstream_data  [ 109] ;
  assign tx_phy_preflop_0 [ 113] = tx_downstream_data  [ 110] ;
  assign tx_phy_preflop_0 [ 114] = tx_downstream_data  [ 111] ;
  assign tx_phy_preflop_0 [ 115] = tx_downstream_data  [ 112] ;
  assign tx_phy_preflop_0 [ 116] = tx_downstream_data  [ 113] ;
  assign tx_phy_preflop_0 [ 117] = tx_downstream_data  [ 114] ;
  assign tx_phy_preflop_0 [ 118] = tx_downstream_data  [ 115] ;
  assign tx_phy_preflop_0 [ 119] = tx_downstream_data  [ 116] ;
  assign tx_phy_preflop_0 [ 120] = tx_downstream_data  [ 117] ;
  assign tx_phy_preflop_0 [ 121] = tx_downstream_data  [ 118] ;
  assign tx_phy_preflop_0 [ 122] = tx_downstream_data  [ 119] ;
  assign tx_phy_preflop_0 [ 123] = tx_downstream_data  [ 120] ;
  assign tx_phy_preflop_0 [ 124] = tx_downstream_data  [ 121] ;
  assign tx_phy_preflop_0 [ 125] = tx_downstream_data  [ 122] ;
  assign tx_phy_preflop_0 [ 126] = tx_downstream_data  [ 123] ;
  assign tx_phy_preflop_0 [ 127] = tx_downstream_data  [ 124] ;
  assign tx_phy_preflop_0 [ 128] = tx_downstream_data  [ 125] ;
  assign tx_phy_preflop_0 [ 129] = tx_downstream_data  [ 126] ;
  assign tx_phy_preflop_0 [ 130] = tx_downstream_data  [ 127] ;
  assign tx_phy_preflop_0 [ 131] = tx_downstream_data  [ 128] ;
  assign tx_phy_preflop_0 [ 132] = tx_downstream_data  [ 129] ;
  assign tx_phy_preflop_0 [ 133] = tx_downstream_data  [ 130] ;
  assign tx_phy_preflop_0 [ 134] = tx_downstream_data  [ 131] ;
  assign tx_phy_preflop_0 [ 135] = tx_downstream_data  [ 132] ;
  assign tx_phy_preflop_0 [ 136] = tx_downstream_data  [ 133] ;
  assign tx_phy_preflop_0 [ 137] = tx_downstream_data  [ 134] ;
  assign tx_phy_preflop_0 [ 138] = tx_downstream_data  [ 135] ;
  assign tx_phy_preflop_0 [ 139] = tx_downstream_data  [ 136] ;
  assign tx_phy_preflop_0 [ 140] = tx_downstream_data  [ 137] ;
  assign tx_phy_preflop_0 [ 141] = tx_downstream_data  [ 138] ;
  assign tx_phy_preflop_0 [ 142] = tx_downstream_data  [ 139] ;
  assign tx_phy_preflop_0 [ 143] = tx_downstream_data  [ 140] ;
  assign tx_phy_preflop_0 [ 144] = tx_downstream_data  [ 141] ;
  assign tx_phy_preflop_0 [ 145] = tx_downstream_data  [ 142] ;
  assign tx_phy_preflop_0 [ 146] = tx_downstream_data  [ 143] ;
  assign tx_phy_preflop_0 [ 147] = tx_downstream_data  [ 144] ;
  assign tx_phy_preflop_0 [ 148] = tx_downstream_data  [ 145] ;
  assign tx_phy_preflop_0 [ 149] = tx_downstream_data  [ 146] ;
  assign tx_phy_preflop_0 [ 150] = tx_downstream_data  [ 147] ;
  assign tx_phy_preflop_0 [ 151] = tx_downstream_data  [ 148] ;
  assign tx_phy_preflop_0 [ 152] = tx_downstream_data  [ 149] ;
  assign tx_phy_preflop_0 [ 153] = tx_downstream_data  [ 150] ;
  assign tx_phy_preflop_0 [ 154] = tx_downstream_data  [ 151] ;
  assign tx_phy_preflop_0 [ 155] = tx_downstream_data  [ 152] ;
  assign tx_phy_preflop_0 [ 156] = tx_downstream_data  [ 153] ;
  assign tx_phy_preflop_0 [ 157] = tx_downstream_data  [ 154] ;
  assign tx_phy_preflop_0 [ 158] = tx_downstream_data  [ 155] ;
  assign tx_phy_preflop_0 [ 159] = tx_downstream_data  [ 156] ;
  assign tx_phy_preflop_1 [   0] = tx_downstream_data  [ 157] ;
  assign tx_phy_preflop_1 [   1] = tx_downstream_data  [ 158] ;
  assign tx_phy_preflop_1 [   2] = tx_downstream_data  [ 159] ;
  assign tx_phy_preflop_1 [   3] = tx_downstream_data  [ 160] ;
  assign tx_phy_preflop_1 [   4] = tx_mrk_userbit[0]          ; // MARKER
  assign tx_phy_preflop_1 [   5] = tx_downstream_data  [ 161] ;
  assign tx_phy_preflop_1 [   6] = tx_downstream_data  [ 162] ;
  assign tx_phy_preflop_1 [   7] = tx_downstream_data  [ 163] ;
  assign tx_phy_preflop_1 [   8] = tx_downstream_data  [ 164] ;
  assign tx_phy_preflop_1 [   9] = tx_downstream_data  [ 165] ;
  assign tx_phy_preflop_1 [  10] = tx_downstream_data  [ 166] ;
  assign tx_phy_preflop_1 [  11] = tx_downstream_data  [ 167] ;
  assign tx_phy_preflop_1 [  12] = tx_downstream_data  [ 168] ;
  assign tx_phy_preflop_1 [  13] = tx_downstream_data  [ 169] ;
  assign tx_phy_preflop_1 [  14] = tx_downstream_data  [ 170] ;
  assign tx_phy_preflop_1 [  15] = tx_downstream_data  [ 171] ;
  assign tx_phy_preflop_1 [  16] = tx_downstream_data  [ 172] ;
  assign tx_phy_preflop_1 [  17] = tx_downstream_data  [ 173] ;
  assign tx_phy_preflop_1 [  18] = tx_downstream_data  [ 174] ;
  assign tx_phy_preflop_1 [  19] = tx_downstream_data  [ 175] ;
  assign tx_phy_preflop_1 [  20] = tx_downstream_data  [ 176] ;
  assign tx_phy_preflop_1 [  21] = tx_downstream_data  [ 177] ;
  assign tx_phy_preflop_1 [  22] = tx_downstream_data  [ 178] ;
  assign tx_phy_preflop_1 [  23] = tx_downstream_data  [ 179] ;
  assign tx_phy_preflop_1 [  24] = tx_downstream_data  [ 180] ;
  assign tx_phy_preflop_1 [  25] = tx_downstream_data  [ 181] ;
  assign tx_phy_preflop_1 [  26] = tx_downstream_data  [ 182] ;
  assign tx_phy_preflop_1 [  27] = tx_downstream_data  [ 183] ;
  assign tx_phy_preflop_1 [  28] = tx_downstream_data  [ 184] ;
  assign tx_phy_preflop_1 [  29] = tx_downstream_data  [ 185] ;
  assign tx_phy_preflop_1 [  30] = tx_downstream_data  [ 186] ;
  assign tx_phy_preflop_1 [  31] = tx_downstream_data  [ 187] ;
  assign tx_phy_preflop_1 [  32] = tx_downstream_data  [ 188] ;
  assign tx_phy_preflop_1 [  33] = tx_downstream_data  [ 189] ;
  assign tx_phy_preflop_1 [  34] = tx_downstream_data  [ 190] ;
  assign tx_phy_preflop_1 [  35] = tx_downstream_data  [ 191] ;
  assign tx_phy_preflop_1 [  36] = tx_downstream_data  [ 192] ;
  assign tx_phy_preflop_1 [  37] = tx_downstream_data  [ 193] ;
  assign tx_phy_preflop_1 [  38] = tx_downstream_data  [ 194] ;
  assign tx_phy_preflop_1 [  39] = tx_downstream_data  [ 195] ;
  assign tx_phy_preflop_1 [  40] = tx_downstream_data  [ 196] ;
  assign tx_phy_preflop_1 [  41] = tx_downstream_data  [ 197] ;
  assign tx_phy_preflop_1 [  42] = tx_downstream_data  [ 198] ;
  assign tx_phy_preflop_1 [  43] = tx_downstream_data  [ 199] ;
  assign tx_phy_preflop_1 [  44] = tx_downstream_data  [ 200] ;
  assign tx_phy_preflop_1 [  45] = tx_downstream_data  [ 201] ;
  assign tx_phy_preflop_1 [  46] = tx_downstream_data  [ 202] ;
  assign tx_phy_preflop_1 [  47] = tx_downstream_data  [ 203] ;
  assign tx_phy_preflop_1 [  48] = tx_downstream_data  [ 204] ;
  assign tx_phy_preflop_1 [  49] = tx_downstream_data  [ 205] ;
  assign tx_phy_preflop_1 [  50] = tx_downstream_data  [ 206] ;
  assign tx_phy_preflop_1 [  51] = tx_downstream_data  [ 207] ;
  assign tx_phy_preflop_1 [  52] = tx_downstream_data  [ 208] ;
  assign tx_phy_preflop_1 [  53] = tx_downstream_data  [ 209] ;
  assign tx_phy_preflop_1 [  54] = tx_downstream_data  [ 210] ;
  assign tx_phy_preflop_1 [  55] = tx_downstream_data  [ 211] ;
  assign tx_phy_preflop_1 [  56] = tx_downstream_data  [ 212] ;
  assign tx_phy_preflop_1 [  57] = tx_downstream_data  [ 213] ;
  assign tx_phy_preflop_1 [  58] = tx_downstream_data  [ 214] ;
  assign tx_phy_preflop_1 [  59] = tx_downstream_data  [ 215] ;
  assign tx_phy_preflop_1 [  60] = tx_downstream_data  [ 216] ;
  assign tx_phy_preflop_1 [  61] = tx_downstream_data  [ 217] ;
  assign tx_phy_preflop_1 [  62] = tx_downstream_data  [ 218] ;
  assign tx_phy_preflop_1 [  63] = tx_downstream_data  [ 219] ;
  assign tx_phy_preflop_1 [  64] = tx_downstream_data  [ 220] ;
  assign tx_phy_preflop_1 [  65] = tx_downstream_data  [ 221] ;
  assign tx_phy_preflop_1 [  66] = tx_downstream_data  [ 222] ;
  assign tx_phy_preflop_1 [  67] = tx_downstream_data  [ 223] ;
  assign tx_phy_preflop_1 [  68] = tx_downstream_data  [ 224] ;
  assign tx_phy_preflop_1 [  69] = tx_downstream_data  [ 225] ;
  assign tx_phy_preflop_1 [  70] = tx_downstream_data  [ 226] ;
  assign tx_phy_preflop_1 [  71] = tx_downstream_data  [ 227] ;
  assign tx_phy_preflop_1 [  72] = tx_downstream_data  [ 228] ;
  assign tx_phy_preflop_1 [  73] = tx_downstream_data  [ 229] ;
  assign tx_phy_preflop_1 [  74] = tx_downstream_data  [ 230] ;
  assign tx_phy_preflop_1 [  75] = tx_downstream_data  [ 231] ;
  assign tx_phy_preflop_1 [  76] = tx_stb_userbit             ; // STROBE
  assign tx_phy_preflop_1 [  77] = tx_downstream_data  [ 232] ;
  assign tx_phy_preflop_1 [  78] = tx_downstream_data  [ 233] ;
  assign tx_phy_preflop_1 [  79] = tx_downstream_data  [ 234] ;
  assign tx_phy_preflop_1 [  80] = tx_downstream_data  [ 235] ;
  assign tx_phy_preflop_1 [  81] = tx_downstream_data  [ 236] ;
  assign tx_phy_preflop_1 [  82] = tx_downstream_data  [ 237] ;
  assign tx_phy_preflop_1 [  83] = tx_downstream_data  [ 238] ;
  assign tx_phy_preflop_1 [  84] = tx_mrk_userbit[1]          ; // MARKER
  assign tx_phy_preflop_1 [  85] = tx_downstream_data  [ 239] ;
  assign tx_phy_preflop_1 [  86] = tx_downstream_data  [ 240] ;
  assign tx_phy_preflop_1 [  87] = tx_downstream_data  [ 241] ;
  assign tx_phy_preflop_1 [  88] = tx_downstream_data  [ 242] ;
  assign tx_phy_preflop_1 [  89] = tx_downstream_data  [ 243] ;
  assign tx_phy_preflop_1 [  90] = tx_downstream_data  [ 244] ;
  assign tx_phy_preflop_1 [  91] = tx_downstream_data  [ 245] ;
  assign tx_phy_preflop_1 [  92] = tx_downstream_data  [ 246] ;
  assign tx_phy_preflop_1 [  93] = tx_downstream_data  [ 247] ;
  assign tx_phy_preflop_1 [  94] = tx_downstream_data  [ 248] ;
  assign tx_phy_preflop_1 [  95] = tx_downstream_data  [ 249] ;
  assign tx_phy_preflop_1 [  96] = tx_downstream_data  [ 250] ;
  assign tx_phy_preflop_1 [  97] = tx_downstream_data  [ 251] ;
  assign tx_phy_preflop_1 [  98] = tx_downstream_data  [ 252] ;
  assign tx_phy_preflop_1 [  99] = tx_downstream_data  [ 253] ;
  assign tx_phy_preflop_1 [ 100] = tx_downstream_data  [ 254] ;
  assign tx_phy_preflop_1 [ 101] = tx_downstream_data  [ 255] ;
  assign tx_phy_preflop_1 [ 102] = tx_downstream_data  [ 256] ;
  assign tx_phy_preflop_1 [ 103] = tx_downstream_data  [ 257] ;
  assign tx_phy_preflop_1 [ 104] = tx_downstream_data  [ 258] ;
  assign tx_phy_preflop_1 [ 105] = tx_downstream_data  [ 259] ;
  assign tx_phy_preflop_1 [ 106] = tx_downstream_data  [ 260] ;
  assign tx_phy_preflop_1 [ 107] = tx_downstream_data  [ 261] ;
  assign tx_phy_preflop_1 [ 108] = tx_downstream_data  [ 262] ;
  assign tx_phy_preflop_1 [ 109] = tx_downstream_data  [ 263] ;
  assign tx_phy_preflop_1 [ 110] = tx_downstream_data  [ 264] ;
  assign tx_phy_preflop_1 [ 111] = tx_downstream_data  [ 265] ;
  assign tx_phy_preflop_1 [ 112] = tx_downstream_data  [ 266] ;
  assign tx_phy_preflop_1 [ 113] = tx_downstream_data  [ 267] ;
  assign tx_phy_preflop_1 [ 114] = tx_downstream_data  [ 268] ;
  assign tx_phy_preflop_1 [ 115] = tx_downstream_data  [ 269] ;
  assign tx_phy_preflop_1 [ 116] = tx_downstream_data  [ 270] ;
  assign tx_phy_preflop_1 [ 117] = tx_downstream_data  [ 271] ;
  assign tx_phy_preflop_1 [ 118] = tx_downstream_data  [ 272] ;
  assign tx_phy_preflop_1 [ 119] = tx_downstream_data  [ 273] ;
  assign tx_phy_preflop_1 [ 120] = tx_downstream_data  [ 274] ;
  assign tx_phy_preflop_1 [ 121] = tx_downstream_data  [ 275] ;
  assign tx_phy_preflop_1 [ 122] = tx_downstream_data  [ 276] ;
  assign tx_phy_preflop_1 [ 123] = tx_downstream_data  [ 277] ;
  assign tx_phy_preflop_1 [ 124] = tx_downstream_data  [ 278] ;
  assign tx_phy_preflop_1 [ 125] = tx_downstream_data  [ 279] ;
  assign tx_phy_preflop_1 [ 126] = tx_downstream_data  [ 280] ;
  assign tx_phy_preflop_1 [ 127] = tx_downstream_data  [ 281] ;
  assign tx_phy_preflop_1 [ 128] = tx_downstream_data  [ 282] ;
  assign tx_phy_preflop_1 [ 129] = tx_downstream_data  [ 283] ;
  assign tx_phy_preflop_1 [ 130] = tx_downstream_data  [ 284] ;
  assign tx_phy_preflop_1 [ 131] = tx_downstream_data  [ 285] ;
  assign tx_phy_preflop_1 [ 132] = tx_downstream_data  [ 286] ;
  assign tx_phy_preflop_1 [ 133] = tx_downstream_data  [ 287] ;
  assign tx_phy_preflop_1 [ 134] = tx_downstream_data  [ 288] ;
  assign tx_phy_preflop_1 [ 135] = tx_downstream_data  [ 289] ;
  assign tx_phy_preflop_1 [ 136] = tx_downstream_data  [ 290] ;
  assign tx_phy_preflop_1 [ 137] = tx_downstream_data  [ 291] ;
  assign tx_phy_preflop_1 [ 138] = tx_downstream_data  [ 292] ;
  assign tx_phy_preflop_1 [ 139] = tx_downstream_data  [ 293] ;
  assign tx_phy_preflop_1 [ 140] = tx_downstream_data  [ 294] ;
  assign tx_phy_preflop_1 [ 141] = tx_downstream_data  [ 295] ;
  assign tx_phy_preflop_1 [ 142] = tx_downstream_data  [ 296] ;
  assign tx_phy_preflop_1 [ 143] = tx_downstream_data  [ 297] ;
  assign tx_phy_preflop_1 [ 144] = tx_downstream_data  [ 298] ;
  assign tx_phy_preflop_1 [ 145] = tx_downstream_data  [ 299] ;
  assign tx_phy_preflop_1 [ 146] = tx_downstream_data  [ 300] ;
  assign tx_phy_preflop_1 [ 147] = tx_downstream_data  [ 301] ;
  assign tx_phy_preflop_1 [ 148] = tx_downstream_data  [ 302] ;
  assign tx_phy_preflop_1 [ 149] = tx_downstream_data  [ 303] ;
  assign tx_phy_preflop_1 [ 150] = tx_downstream_data  [ 304] ;
  assign tx_phy_preflop_1 [ 151] = tx_downstream_data  [ 305] ;
  assign tx_phy_preflop_1 [ 152] = tx_downstream_data  [ 306] ;
  assign tx_phy_preflop_1 [ 153] = tx_downstream_data  [ 307] ;
  assign tx_phy_preflop_1 [ 154] = tx_downstream_data  [ 308] ;
  assign tx_phy_preflop_1 [ 155] = tx_downstream_data  [ 309] ;
  assign tx_phy_preflop_1 [ 156] = tx_downstream_data  [ 310] ;
  assign tx_phy_preflop_1 [ 157] = tx_downstream_data  [ 311] ;
  assign tx_phy_preflop_1 [ 158] = tx_downstream_data  [ 312] ;
  assign tx_phy_preflop_1 [ 159] = tx_downstream_data  [ 313] ;
  assign tx_phy_preflop_2 [   0] = tx_downstream_data  [ 314] ;
  assign tx_phy_preflop_2 [   1] = tx_downstream_data  [ 315] ;
  assign tx_phy_preflop_2 [   2] = tx_downstream_data  [ 316] ;
  assign tx_phy_preflop_2 [   3] = tx_downstream_data  [ 317] ;
  assign tx_phy_preflop_2 [   4] = tx_mrk_userbit[0]          ; // MARKER
  assign tx_phy_preflop_2 [   5] = tx_downstream_data  [ 318] ;
  assign tx_phy_preflop_2 [   6] = tx_downstream_data  [ 319] ;
  assign tx_phy_preflop_2 [   7] = tx_downstream_data  [ 320] ;
  assign tx_phy_preflop_2 [   8] = tx_downstream_data  [ 321] ;
  assign tx_phy_preflop_2 [   9] = tx_downstream_data  [ 322] ;
  assign tx_phy_preflop_2 [  10] = tx_downstream_data  [ 323] ;
  assign tx_phy_preflop_2 [  11] = tx_downstream_data  [ 324] ;
  assign tx_phy_preflop_2 [  12] = tx_downstream_data  [ 325] ;
  assign tx_phy_preflop_2 [  13] = tx_downstream_data  [ 326] ;
  assign tx_phy_preflop_2 [  14] = tx_downstream_data  [ 327] ;
  assign tx_phy_preflop_2 [  15] = tx_downstream_data  [ 328] ;
  assign tx_phy_preflop_2 [  16] = tx_downstream_data  [ 329] ;
  assign tx_phy_preflop_2 [  17] = tx_downstream_data  [ 330] ;
  assign tx_phy_preflop_2 [  18] = tx_downstream_data  [ 331] ;
  assign tx_phy_preflop_2 [  19] = tx_downstream_data  [ 332] ;
  assign tx_phy_preflop_2 [  20] = tx_downstream_data  [ 333] ;
  assign tx_phy_preflop_2 [  21] = tx_downstream_data  [ 334] ;
  assign tx_phy_preflop_2 [  22] = tx_downstream_data  [ 335] ;
  assign tx_phy_preflop_2 [  23] = tx_downstream_data  [ 336] ;
  assign tx_phy_preflop_2 [  24] = tx_downstream_data  [ 337] ;
  assign tx_phy_preflop_2 [  25] = tx_downstream_data  [ 338] ;
  assign tx_phy_preflop_2 [  26] = tx_downstream_data  [ 339] ;
  assign tx_phy_preflop_2 [  27] = tx_downstream_data  [ 340] ;
  assign tx_phy_preflop_2 [  28] = tx_downstream_data  [ 341] ;
  assign tx_phy_preflop_2 [  29] = tx_downstream_data  [ 342] ;
  assign tx_phy_preflop_2 [  30] = tx_downstream_data  [ 343] ;
  assign tx_phy_preflop_2 [  31] = tx_downstream_data  [ 344] ;
  assign tx_phy_preflop_2 [  32] = tx_downstream_data  [ 345] ;
  assign tx_phy_preflop_2 [  33] = tx_downstream_data  [ 346] ;
  assign tx_phy_preflop_2 [  34] = tx_downstream_data  [ 347] ;
  assign tx_phy_preflop_2 [  35] = tx_downstream_data  [ 348] ;
  assign tx_phy_preflop_2 [  36] = tx_downstream_data  [ 349] ;
  assign tx_phy_preflop_2 [  37] = tx_downstream_data  [ 350] ;
  assign tx_phy_preflop_2 [  38] = tx_downstream_data  [ 351] ;
  assign tx_phy_preflop_2 [  39] = tx_downstream_data  [ 352] ;
  assign tx_phy_preflop_2 [  40] = tx_downstream_data  [ 353] ;
  assign tx_phy_preflop_2 [  41] = tx_downstream_data  [ 354] ;
  assign tx_phy_preflop_2 [  42] = tx_downstream_data  [ 355] ;
  assign tx_phy_preflop_2 [  43] = tx_downstream_data  [ 356] ;
  assign tx_phy_preflop_2 [  44] = tx_downstream_data  [ 357] ;
  assign tx_phy_preflop_2 [  45] = tx_downstream_data  [ 358] ;
  assign tx_phy_preflop_2 [  46] = tx_downstream_data  [ 359] ;
  assign tx_phy_preflop_2 [  47] = tx_downstream_data  [ 360] ;
  assign tx_phy_preflop_2 [  48] = tx_downstream_data  [ 361] ;
  assign tx_phy_preflop_2 [  49] = tx_downstream_data  [ 362] ;
  assign tx_phy_preflop_2 [  50] = tx_downstream_data  [ 363] ;
  assign tx_phy_preflop_2 [  51] = tx_downstream_data  [ 364] ;
  assign tx_phy_preflop_2 [  52] = tx_downstream_data  [ 365] ;
  assign tx_phy_preflop_2 [  53] = tx_downstream_data  [ 366] ;
  assign tx_phy_preflop_2 [  54] = tx_downstream_data  [ 367] ;
  assign tx_phy_preflop_2 [  55] = tx_downstream_data  [ 368] ;
  assign tx_phy_preflop_2 [  56] = tx_downstream_data  [ 369] ;
  assign tx_phy_preflop_2 [  57] = tx_downstream_data  [ 370] ;
  assign tx_phy_preflop_2 [  58] = tx_downstream_data  [ 371] ;
  assign tx_phy_preflop_2 [  59] = tx_downstream_data  [ 372] ;
  assign tx_phy_preflop_2 [  60] = tx_downstream_data  [ 373] ;
  assign tx_phy_preflop_2 [  61] = tx_downstream_data  [ 374] ;
  assign tx_phy_preflop_2 [  62] = tx_downstream_data  [ 375] ;
  assign tx_phy_preflop_2 [  63] = tx_downstream_data  [ 376] ;
  assign tx_phy_preflop_2 [  64] = tx_downstream_data  [ 377] ;
  assign tx_phy_preflop_2 [  65] = tx_downstream_data  [ 378] ;
  assign tx_phy_preflop_2 [  66] = tx_downstream_data  [ 379] ;
  assign tx_phy_preflop_2 [  67] = tx_downstream_data  [ 380] ;
  assign tx_phy_preflop_2 [  68] = tx_downstream_data  [ 381] ;
  assign tx_phy_preflop_2 [  69] = tx_downstream_data  [ 382] ;
  assign tx_phy_preflop_2 [  70] = tx_downstream_data  [ 383] ;
  assign tx_phy_preflop_2 [  71] = tx_downstream_data  [ 384] ;
  assign tx_phy_preflop_2 [  72] = tx_downstream_data  [ 385] ;
  assign tx_phy_preflop_2 [  73] = tx_downstream_data  [ 386] ;
  assign tx_phy_preflop_2 [  74] = tx_downstream_data  [ 387] ;
  assign tx_phy_preflop_2 [  75] = tx_downstream_data  [ 388] ;
  assign tx_phy_preflop_2 [  76] = tx_stb_userbit             ; // STROBE
  assign tx_phy_preflop_2 [  77] = tx_downstream_data  [ 389] ;
  assign tx_phy_preflop_2 [  78] = tx_downstream_data  [ 390] ;
  assign tx_phy_preflop_2 [  79] = tx_downstream_data  [ 391] ;
  assign tx_phy_preflop_2 [  80] = tx_downstream_data  [ 392] ;
  assign tx_phy_preflop_2 [  81] = tx_downstream_data  [ 393] ;
  assign tx_phy_preflop_2 [  82] = tx_downstream_data  [ 394] ;
  assign tx_phy_preflop_2 [  83] = tx_downstream_data  [ 395] ;
  assign tx_phy_preflop_2 [  84] = tx_mrk_userbit[1]          ; // MARKER
  assign tx_phy_preflop_2 [  85] = tx_downstream_data  [ 396] ;
  assign tx_phy_preflop_2 [  86] = tx_downstream_data  [ 397] ;
  assign tx_phy_preflop_2 [  87] = tx_downstream_data  [ 398] ;
  assign tx_phy_preflop_2 [  88] = tx_downstream_data  [ 399] ;
  assign tx_phy_preflop_2 [  89] = tx_downstream_data  [ 400] ;
  assign tx_phy_preflop_2 [  90] = tx_downstream_data  [ 401] ;
  assign tx_phy_preflop_2 [  91] = tx_downstream_data  [ 402] ;
  assign tx_phy_preflop_2 [  92] = tx_downstream_data  [ 403] ;
  assign tx_phy_preflop_2 [  93] = tx_downstream_data  [ 404] ;
  assign tx_phy_preflop_2 [  94] = tx_downstream_data  [ 405] ;
  assign tx_phy_preflop_2 [  95] = tx_downstream_data  [ 406] ;
  assign tx_phy_preflop_2 [  96] = tx_downstream_data  [ 407] ;
  assign tx_phy_preflop_2 [  97] = tx_downstream_data  [ 408] ;
  assign tx_phy_preflop_2 [  98] = tx_downstream_data  [ 409] ;
  assign tx_phy_preflop_2 [  99] = tx_downstream_data  [ 410] ;
  assign tx_phy_preflop_2 [ 100] = tx_downstream_data  [ 411] ;
  assign tx_phy_preflop_2 [ 101] = tx_downstream_data  [ 412] ;
  assign tx_phy_preflop_2 [ 102] = tx_downstream_data  [ 413] ;
  assign tx_phy_preflop_2 [ 103] = tx_downstream_data  [ 414] ;
  assign tx_phy_preflop_2 [ 104] = tx_downstream_data  [ 415] ;
  assign tx_phy_preflop_2 [ 105] = tx_downstream_data  [ 416] ;
  assign tx_phy_preflop_2 [ 106] = tx_downstream_data  [ 417] ;
  assign tx_phy_preflop_2 [ 107] = tx_downstream_data  [ 418] ;
  assign tx_phy_preflop_2 [ 108] = tx_downstream_data  [ 419] ;
  assign tx_phy_preflop_2 [ 109] = tx_downstream_data  [ 420] ;
  assign tx_phy_preflop_2 [ 110] = tx_downstream_data  [ 421] ;
  assign tx_phy_preflop_2 [ 111] = tx_downstream_data  [ 422] ;
  assign tx_phy_preflop_2 [ 112] = tx_downstream_data  [ 423] ;
  assign tx_phy_preflop_2 [ 113] = tx_downstream_data  [ 424] ;
  assign tx_phy_preflop_2 [ 114] = tx_downstream_data  [ 425] ;
  assign tx_phy_preflop_2 [ 115] = tx_downstream_data  [ 426] ;
  assign tx_phy_preflop_2 [ 116] = tx_downstream_data  [ 427] ;
  assign tx_phy_preflop_2 [ 117] = tx_downstream_data  [ 428] ;
  assign tx_phy_preflop_2 [ 118] = tx_downstream_data  [ 429] ;
  assign tx_phy_preflop_2 [ 119] = tx_downstream_data  [ 430] ;
  assign tx_phy_preflop_2 [ 120] = tx_downstream_data  [ 431] ;
  assign tx_phy_preflop_2 [ 121] = tx_downstream_data  [ 432] ;
  assign tx_phy_preflop_2 [ 122] = tx_downstream_data  [ 433] ;
  assign tx_phy_preflop_2 [ 123] = tx_downstream_data  [ 434] ;
  assign tx_phy_preflop_2 [ 124] = tx_downstream_data  [ 435] ;
  assign tx_phy_preflop_2 [ 125] = tx_downstream_data  [ 436] ;
  assign tx_phy_preflop_2 [ 126] = tx_downstream_data  [ 437] ;
  assign tx_phy_preflop_2 [ 127] = tx_downstream_data  [ 438] ;
  assign tx_phy_preflop_2 [ 128] = tx_downstream_data  [ 439] ;
  assign tx_phy_preflop_2 [ 129] = tx_downstream_data  [ 440] ;
  assign tx_phy_preflop_2 [ 130] = tx_downstream_data  [ 441] ;
  assign tx_phy_preflop_2 [ 131] = tx_downstream_data  [ 442] ;
  assign tx_phy_preflop_2 [ 132] = tx_downstream_data  [ 443] ;
  assign tx_phy_preflop_2 [ 133] = tx_downstream_data  [ 444] ;
  assign tx_phy_preflop_2 [ 134] = tx_downstream_data  [ 445] ;
  assign tx_phy_preflop_2 [ 135] = tx_downstream_data  [ 446] ;
  assign tx_phy_preflop_2 [ 136] = tx_downstream_data  [ 447] ;
  assign tx_phy_preflop_2 [ 137] = tx_downstream_data  [ 448] ;
  assign tx_phy_preflop_2 [ 138] = tx_downstream_data  [ 449] ;
  assign tx_phy_preflop_2 [ 139] = tx_downstream_data  [ 450] ;
  assign tx_phy_preflop_2 [ 140] = tx_downstream_data  [ 451] ;
  assign tx_phy_preflop_2 [ 141] = tx_downstream_data  [ 452] ;
  assign tx_phy_preflop_2 [ 142] = tx_downstream_data  [ 453] ;
  assign tx_phy_preflop_2 [ 143] = tx_downstream_data  [ 454] ;
  assign tx_phy_preflop_2 [ 144] = tx_downstream_data  [ 455] ;
  assign tx_phy_preflop_2 [ 145] = tx_downstream_data  [ 456] ;
  assign tx_phy_preflop_2 [ 146] = tx_downstream_data  [ 457] ;
  assign tx_phy_preflop_2 [ 147] = tx_downstream_data  [ 458] ;
  assign tx_phy_preflop_2 [ 148] = tx_downstream_data  [ 459] ;
  assign tx_phy_preflop_2 [ 149] = tx_downstream_data  [ 460] ;
  assign tx_phy_preflop_2 [ 150] = tx_downstream_data  [ 461] ;
  assign tx_phy_preflop_2 [ 151] = tx_downstream_data  [ 462] ;
  assign tx_phy_preflop_2 [ 152] = tx_downstream_data  [ 463] ;
  assign tx_phy_preflop_2 [ 153] = tx_downstream_data  [ 464] ;
  assign tx_phy_preflop_2 [ 154] = tx_downstream_data  [ 465] ;
  assign tx_phy_preflop_2 [ 155] = tx_downstream_data  [ 466] ;
  assign tx_phy_preflop_2 [ 156] = tx_downstream_data  [ 467] ;
  assign tx_phy_preflop_2 [ 157] = tx_downstream_data  [ 468] ;
  assign tx_phy_preflop_2 [ 158] = tx_downstream_data  [ 469] ;
  assign tx_phy_preflop_2 [ 159] = tx_downstream_data  [ 470] ;
  assign tx_phy_preflop_3 [   0] = tx_downstream_data  [ 471] ;
  assign tx_phy_preflop_3 [   1] = tx_downstream_data  [ 472] ;
  assign tx_phy_preflop_3 [   2] = tx_downstream_data  [ 473] ;
  assign tx_phy_preflop_3 [   3] = tx_downstream_data  [ 474] ;
  assign tx_phy_preflop_3 [   4] = tx_mrk_userbit[0]          ; // MARKER
  assign tx_phy_preflop_3 [   5] = tx_downstream_data  [ 475] ;
  assign tx_phy_preflop_3 [   6] = tx_downstream_data  [ 476] ;
  assign tx_phy_preflop_3 [   7] = tx_downstream_data  [ 477] ;
  assign tx_phy_preflop_3 [   8] = tx_downstream_data  [ 478] ;
  assign tx_phy_preflop_3 [   9] = tx_downstream_data  [ 479] ;
  assign tx_phy_preflop_3 [  10] = tx_downstream_data  [ 480] ;
  assign tx_phy_preflop_3 [  11] = tx_downstream_data  [ 481] ;
  assign tx_phy_preflop_3 [  12] = tx_downstream_data  [ 482] ;
  assign tx_phy_preflop_3 [  13] = tx_downstream_data  [ 483] ;
  assign tx_phy_preflop_3 [  14] = tx_downstream_data  [ 484] ;
  assign tx_phy_preflop_3 [  15] = tx_downstream_data  [ 485] ;
  assign tx_phy_preflop_3 [  16] = tx_downstream_data  [ 486] ;
  assign tx_phy_preflop_3 [  17] = tx_downstream_data  [ 487] ;
  assign tx_phy_preflop_3 [  18] = tx_downstream_data  [ 488] ;
  assign tx_phy_preflop_3 [  19] = tx_downstream_data  [ 489] ;
  assign tx_phy_preflop_3 [  20] = tx_downstream_data  [ 490] ;
  assign tx_phy_preflop_3 [  21] = tx_downstream_data  [ 491] ;
  assign tx_phy_preflop_3 [  22] = tx_downstream_data  [ 492] ;
  assign tx_phy_preflop_3 [  23] = tx_downstream_data  [ 493] ;
  assign tx_phy_preflop_3 [  24] = tx_downstream_data  [ 494] ;
  assign tx_phy_preflop_3 [  25] = tx_downstream_data  [ 495] ;
  assign tx_phy_preflop_3 [  26] = tx_downstream_data  [ 496] ;
  assign tx_phy_preflop_3 [  27] = tx_downstream_data  [ 497] ;
  assign tx_phy_preflop_3 [  28] = tx_downstream_data  [ 498] ;
  assign tx_phy_preflop_3 [  29] = tx_downstream_data  [ 499] ;
  assign tx_phy_preflop_3 [  30] = tx_downstream_data  [ 500] ;
  assign tx_phy_preflop_3 [  31] = tx_downstream_data  [ 501] ;
  assign tx_phy_preflop_3 [  32] = tx_downstream_data  [ 502] ;
  assign tx_phy_preflop_3 [  33] = tx_downstream_data  [ 503] ;
  assign tx_phy_preflop_3 [  34] = tx_downstream_data  [ 504] ;
  assign tx_phy_preflop_3 [  35] = tx_downstream_data  [ 505] ;
  assign tx_phy_preflop_3 [  36] = tx_downstream_data  [ 506] ;
  assign tx_phy_preflop_3 [  37] = tx_downstream_data  [ 507] ;
  assign tx_phy_preflop_3 [  38] = tx_downstream_data  [ 508] ;
  assign tx_phy_preflop_3 [  39] = tx_downstream_data  [ 509] ;
  assign tx_phy_preflop_3 [  40] = tx_downstream_data  [ 510] ;
  assign tx_phy_preflop_3 [  41] = tx_downstream_data  [ 511] ;
  assign tx_phy_preflop_3 [  42] = tx_downstream_data  [ 512] ;
  assign tx_phy_preflop_3 [  43] = tx_downstream_data  [ 513] ;
  assign tx_phy_preflop_3 [  44] = tx_downstream_data  [ 514] ;
  assign tx_phy_preflop_3 [  45] = tx_downstream_data  [ 515] ;
  assign tx_phy_preflop_3 [  46] = tx_downstream_data  [ 516] ;
  assign tx_phy_preflop_3 [  47] = tx_downstream_data  [ 517] ;
  assign tx_phy_preflop_3 [  48] = tx_downstream_data  [ 518] ;
  assign tx_phy_preflop_3 [  49] = tx_downstream_data  [ 519] ;
  assign tx_phy_preflop_3 [  50] = tx_downstream_data  [ 520] ;
  assign tx_phy_preflop_3 [  51] = tx_downstream_data  [ 521] ;
  assign tx_phy_preflop_3 [  52] = tx_downstream_data  [ 522] ;
  assign tx_phy_preflop_3 [  53] = tx_downstream_data  [ 523] ;
  assign tx_phy_preflop_3 [  54] = tx_downstream_data  [ 524] ;
  assign tx_phy_preflop_3 [  55] = tx_downstream_data  [ 525] ;
  assign tx_phy_preflop_3 [  56] = tx_downstream_data  [ 526] ;
  assign tx_phy_preflop_3 [  57] = tx_downstream_data  [ 527] ;
  assign tx_phy_preflop_3 [  58] = tx_downstream_data  [ 528] ;
  assign tx_phy_preflop_3 [  59] = tx_downstream_data  [ 529] ;
  assign tx_phy_preflop_3 [  60] = tx_downstream_data  [ 530] ;
  assign tx_phy_preflop_3 [  61] = tx_downstream_data  [ 531] ;
  assign tx_phy_preflop_3 [  62] = tx_downstream_data  [ 532] ;
  assign tx_phy_preflop_3 [  63] = tx_downstream_data  [ 533] ;
  assign tx_phy_preflop_3 [  64] = tx_downstream_data  [ 534] ;
  assign tx_phy_preflop_3 [  65] = tx_downstream_data  [ 535] ;
  assign tx_phy_preflop_3 [  66] = tx_downstream_data  [ 536] ;
  assign tx_phy_preflop_3 [  67] = tx_downstream_data  [ 537] ;
  assign tx_phy_preflop_3 [  68] = tx_downstream_data  [ 538] ;
  assign tx_phy_preflop_3 [  69] = tx_downstream_data  [ 539] ;
  assign tx_phy_preflop_3 [  70] = tx_downstream_data  [ 540] ;
  assign tx_phy_preflop_3 [  71] = tx_downstream_data  [ 541] ;
  assign tx_phy_preflop_3 [  72] = tx_downstream_data  [ 542] ;
  assign tx_phy_preflop_3 [  73] = tx_downstream_data  [ 543] ;
  assign tx_phy_preflop_3 [  74] = tx_downstream_data  [ 544] ;
  assign tx_phy_preflop_3 [  75] = tx_downstream_data  [ 545] ;
  assign tx_phy_preflop_3 [  76] = tx_stb_userbit             ; // STROBE
  assign tx_phy_preflop_3 [  77] = tx_downstream_data  [ 546] ;
  assign tx_phy_preflop_3 [  78] = tx_downstream_data  [ 547] ;
  assign tx_phy_preflop_3 [  79] = tx_downstream_data  [ 548] ;
  assign tx_phy_preflop_3 [  80] = tx_downstream_data  [ 549] ;
  assign tx_phy_preflop_3 [  81] = tx_downstream_data  [ 550] ;
  assign tx_phy_preflop_3 [  82] = tx_downstream_data  [ 551] ;
  assign tx_phy_preflop_3 [  83] = tx_downstream_data  [ 552] ;
  assign tx_phy_preflop_3 [  84] = tx_mrk_userbit[1]          ; // MARKER
  assign tx_phy_preflop_3 [  85] = tx_downstream_data  [ 553] ;
  assign tx_phy_preflop_3 [  86] = tx_downstream_data  [ 554] ;
  assign tx_phy_preflop_3 [  87] = tx_downstream_data  [ 555] ;
  assign tx_phy_preflop_3 [  88] = tx_downstream_data  [ 556] ;
  assign tx_phy_preflop_3 [  89] = tx_downstream_data  [ 557] ;
  assign tx_phy_preflop_3 [  90] = tx_downstream_data  [ 558] ;
  assign tx_phy_preflop_3 [  91] = tx_downstream_data  [ 559] ;
  assign tx_phy_preflop_3 [  92] = tx_downstream_data  [ 560] ;
  assign tx_phy_preflop_3 [  93] = tx_downstream_data  [ 561] ;
  assign tx_phy_preflop_3 [  94] = tx_downstream_data  [ 562] ;
  assign tx_phy_preflop_3 [  95] = tx_downstream_data  [ 563] ;
  assign tx_phy_preflop_3 [  96] = tx_downstream_data  [ 564] ;
  assign tx_phy_preflop_3 [  97] = tx_downstream_data  [ 565] ;
  assign tx_phy_preflop_3 [  98] = tx_downstream_data  [ 566] ;
  assign tx_phy_preflop_3 [  99] = tx_downstream_data  [ 567] ;
  assign tx_phy_preflop_3 [ 100] = tx_downstream_data  [ 568] ;
  assign tx_phy_preflop_3 [ 101] = tx_downstream_data  [ 569] ;
  assign tx_phy_preflop_3 [ 102] = tx_downstream_data  [ 570] ;
  assign tx_phy_preflop_3 [ 103] = tx_downstream_data  [ 571] ;
  assign tx_phy_preflop_3 [ 104] = tx_downstream_data  [ 572] ;
  assign tx_phy_preflop_3 [ 105] = tx_downstream_data  [ 573] ;
  assign tx_phy_preflop_3 [ 106] = tx_downstream_data  [ 574] ;
  assign tx_phy_preflop_3 [ 107] = tx_downstream_data  [ 575] ;
  assign tx_phy_preflop_3 [ 108] = tx_downstream_data  [ 576] ;
  assign tx_phy_preflop_3 [ 109] = tx_downstream_data  [ 577] ;
  assign tx_phy_preflop_3 [ 110] = tx_downstream_data  [ 578] ;
  assign tx_phy_preflop_3 [ 111] = tx_downstream_data  [ 579] ;
  assign tx_phy_preflop_3 [ 112] = tx_downstream_data  [ 580] ;
  assign tx_phy_preflop_3 [ 113] = tx_downstream_data  [ 581] ;
  assign tx_phy_preflop_3 [ 114] = tx_downstream_data  [ 582] ;
  assign tx_phy_preflop_3 [ 115] = tx_downstream_data  [ 583] ;
  assign tx_phy_preflop_3 [ 116] = tx_downstream_data  [ 584] ;
  assign tx_phy_preflop_3 [ 117] = tx_downstream_data  [ 585] ;
  assign tx_phy_preflop_3 [ 118] = tx_downstream_data  [ 586] ;
  assign tx_phy_preflop_3 [ 119] = tx_downstream_data  [ 587] ;
  assign tx_phy_preflop_3 [ 120] = tx_downstream_data  [ 588] ;
  assign tx_phy_preflop_3 [ 121] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 122] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 123] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 124] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 125] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 126] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 127] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 128] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 129] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 130] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 131] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 132] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 133] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 134] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 135] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 136] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 137] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 138] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 139] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 140] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 141] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 142] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 143] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 144] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 145] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 146] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 147] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 148] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 149] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 150] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 151] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 152] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 153] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 154] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 155] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 156] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 157] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 158] = 1'b0                       ;
  assign tx_phy_preflop_3 [ 159] = 1'b0                       ;
// TX Section
//////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////
// RX Section

//   RX_CH_WIDTH           = 160; // Gen2 running at Half Rate
//   RX_DATA_WIDTH         = 157; // Usable Data per Channel
//   RX_PERSISTENT_STROBE  = 1'b1;
//   RX_PERSISTENT_MARKER  = 1'b1;
//   RX_STROBE_GEN2_LOC    = 'd76;
//   RX_MARKER_GEN2_LOC    = 'd4;
//   RX_STROBE_GEN1_LOC    = 'd38;
//   RX_MARKER_GEN1_LOC    = 'd39;
//   RX_ENABLE_STROBE      = 1'b1;
//   RX_ENABLE_MARKER      = 1'b1;
//   RX_DBI_PRESENT        = 1'b0;
//   RX_REG_PHY            = 1'b0;

  localparam RX_REG_PHY    = 1'b0;  // If set, this enables boundary FF for timing reasons

  logic [ 159:   0]                              rx_phy_postflop_0             ;
  logic [ 159:   0]                              rx_phy_postflop_1             ;
  logic [ 159:   0]                              rx_phy_postflop_2             ;
  logic [ 159:   0]                              rx_phy_postflop_3             ;
  logic [ 159:   0]                              rx_phy_flop_0_reg             ;
  logic [ 159:   0]                              rx_phy_flop_1_reg             ;
  logic [ 159:   0]                              rx_phy_flop_2_reg             ;
  logic [ 159:   0]                              rx_phy_flop_3_reg             ;

  always_ff @(posedge clk_rd or negedge rst_rd_n)
  if (~rst_rd_n)
  begin
    rx_phy_flop_0_reg                       <= 160'b0                                  ;
    rx_phy_flop_1_reg                       <= 160'b0                                  ;
    rx_phy_flop_2_reg                       <= 160'b0                                  ;
    rx_phy_flop_3_reg                       <= 160'b0                                  ;
  end
  else
  begin
    rx_phy_flop_0_reg                       <= rx_phy0                                 ;
    rx_phy_flop_1_reg                       <= rx_phy1                                 ;
    rx_phy_flop_2_reg                       <= rx_phy2                                 ;
    rx_phy_flop_3_reg                       <= rx_phy3                                 ;
  end


  assign rx_phy_postflop_0                  = RX_REG_PHY ? rx_phy_flop_0_reg : rx_phy0               ;
  assign rx_phy_postflop_1                  = RX_REG_PHY ? rx_phy_flop_1_reg : rx_phy1               ;
  assign rx_phy_postflop_2                  = RX_REG_PHY ? rx_phy_flop_2_reg : rx_phy2               ;
  assign rx_phy_postflop_3                  = RX_REG_PHY ? rx_phy_flop_3_reg : rx_phy3               ;

  assign rx_upstream_data    [   0] = rx_phy_postflop_0 [   0];
  assign rx_upstream_data    [   1] = rx_phy_postflop_0 [   1];
  assign rx_upstream_data    [   2] = rx_phy_postflop_0 [   2];
  assign rx_upstream_data    [   3] = rx_phy_postflop_0 [   3];
//       MARKER                     = rx_phy_postflop_0 [   4]
  assign rx_upstream_data    [   4] = rx_phy_postflop_0 [   5];
  assign rx_upstream_data    [   5] = rx_phy_postflop_0 [   6];
  assign rx_upstream_data    [   6] = rx_phy_postflop_0 [   7];
  assign rx_upstream_data    [   7] = rx_phy_postflop_0 [   8];
  assign rx_upstream_data    [   8] = rx_phy_postflop_0 [   9];
  assign rx_upstream_data    [   9] = rx_phy_postflop_0 [  10];
  assign rx_upstream_data    [  10] = rx_phy_postflop_0 [  11];
  assign rx_upstream_data    [  11] = rx_phy_postflop_0 [  12];
  assign rx_upstream_data    [  12] = rx_phy_postflop_0 [  13];
  assign rx_upstream_data    [  13] = rx_phy_postflop_0 [  14];
  assign rx_upstream_data    [  14] = rx_phy_postflop_0 [  15];
  assign rx_upstream_data    [  15] = rx_phy_postflop_0 [  16];
  assign rx_upstream_data    [  16] = rx_phy_postflop_0 [  17];
  assign rx_upstream_data    [  17] = rx_phy_postflop_0 [  18];
  assign rx_upstream_data    [  18] = rx_phy_postflop_0 [  19];
  assign rx_upstream_data    [  19] = rx_phy_postflop_0 [  20];
  assign rx_upstream_data    [  20] = rx_phy_postflop_0 [  21];
  assign rx_upstream_data    [  21] = rx_phy_postflop_0 [  22];
  assign rx_upstream_data    [  22] = rx_phy_postflop_0 [  23];
  assign rx_upstream_data    [  23] = rx_phy_postflop_0 [  24];
  assign rx_upstream_data    [  24] = rx_phy_postflop_0 [  25];
  assign rx_upstream_data    [  25] = rx_phy_postflop_0 [  26];
  assign rx_upstream_data    [  26] = rx_phy_postflop_0 [  27];
  assign rx_upstream_data    [  27] = rx_phy_postflop_0 [  28];
  assign rx_upstream_data    [  28] = rx_phy_postflop_0 [  29];
  assign rx_upstream_data    [  29] = rx_phy_postflop_0 [  30];
  assign rx_upstream_data    [  30] = rx_phy_postflop_0 [  31];
  assign rx_upstream_data    [  31] = rx_phy_postflop_0 [  32];
  assign rx_upstream_data    [  32] = rx_phy_postflop_0 [  33];
  assign rx_upstream_data    [  33] = rx_phy_postflop_0 [  34];
  assign rx_upstream_data    [  34] = rx_phy_postflop_0 [  35];
  assign rx_upstream_data    [  35] = rx_phy_postflop_0 [  36];
  assign rx_upstream_data    [  36] = rx_phy_postflop_0 [  37];
  assign rx_upstream_data    [  37] = rx_phy_postflop_0 [  38];
  assign rx_upstream_data    [  38] = rx_phy_postflop_0 [  39];
  assign rx_upstream_data    [  39] = rx_phy_postflop_0 [  40];
  assign rx_upstream_data    [  40] = rx_phy_postflop_0 [  41];
  assign rx_upstream_data    [  41] = rx_phy_postflop_0 [  42];
  assign rx_upstream_data    [  42] = rx_phy_postflop_0 [  43];
  assign rx_upstream_data    [  43] = rx_phy_postflop_0 [  44];
  assign rx_upstream_data    [  44] = rx_phy_postflop_0 [  45];
  assign rx_upstream_data    [  45] = rx_phy_postflop_0 [  46];
  assign rx_upstream_data    [  46] = rx_phy_postflop_0 [  47];
  assign rx_upstream_data    [  47] = rx_phy_postflop_0 [  48];
  assign rx_upstream_data    [  48] = rx_phy_postflop_0 [  49];
  assign rx_upstream_data    [  49] = rx_phy_postflop_0 [  50];
  assign rx_upstream_data    [  50] = rx_phy_postflop_0 [  51];
  assign rx_upstream_data    [  51] = rx_phy_postflop_0 [  52];
  assign rx_upstream_data    [  52] = rx_phy_postflop_0 [  53];
  assign rx_upstream_data    [  53] = rx_phy_postflop_0 [  54];
  assign rx_upstream_data    [  54] = rx_phy_postflop_0 [  55];
  assign rx_upstream_data    [  55] = rx_phy_postflop_0 [  56];
  assign rx_upstream_data    [  56] = rx_phy_postflop_0 [  57];
  assign rx_upstream_data    [  57] = rx_phy_postflop_0 [  58];
  assign rx_upstream_data    [  58] = rx_phy_postflop_0 [  59];
  assign rx_upstream_data    [  59] = rx_phy_postflop_0 [  60];
  assign rx_upstream_data    [  60] = rx_phy_postflop_0 [  61];
  assign rx_upstream_data    [  61] = rx_phy_postflop_0 [  62];
  assign rx_upstream_data    [  62] = rx_phy_postflop_0 [  63];
  assign rx_upstream_data    [  63] = rx_phy_postflop_0 [  64];
  assign rx_upstream_data    [  64] = rx_phy_postflop_0 [  65];
  assign rx_upstream_data    [  65] = rx_phy_postflop_0 [  66];
  assign rx_upstream_data    [  66] = rx_phy_postflop_0 [  67];
  assign rx_upstream_data    [  67] = rx_phy_postflop_0 [  68];
  assign rx_upstream_data    [  68] = rx_phy_postflop_0 [  69];
  assign rx_upstream_data    [  69] = rx_phy_postflop_0 [  70];
  assign rx_upstream_data    [  70] = rx_phy_postflop_0 [  71];
  assign rx_upstream_data    [  71] = rx_phy_postflop_0 [  72];
  assign rx_upstream_data    [  72] = rx_phy_postflop_0 [  73];
  assign rx_upstream_data    [  73] = rx_phy_postflop_0 [  74];
  assign rx_upstream_data    [  74] = rx_phy_postflop_0 [  75];
//       STROBE                     = rx_phy_postflop_0 [  76]
  assign rx_upstream_data    [  75] = rx_phy_postflop_0 [  77];
  assign rx_upstream_data    [  76] = rx_phy_postflop_0 [  78];
  assign rx_upstream_data    [  77] = rx_phy_postflop_0 [  79];
  assign rx_upstream_data    [  78] = rx_phy_postflop_0 [  80];
  assign rx_upstream_data    [  79] = rx_phy_postflop_0 [  81];
  assign rx_upstream_data    [  80] = rx_phy_postflop_0 [  82];
  assign rx_upstream_data    [  81] = rx_phy_postflop_0 [  83];
//       MARKER                     = rx_phy_postflop_0 [  84]
  assign rx_upstream_data    [  82] = rx_phy_postflop_0 [  85];
  assign rx_upstream_data    [  83] = rx_phy_postflop_0 [  86];
  assign rx_upstream_data    [  84] = rx_phy_postflop_0 [  87];
  assign rx_upstream_data    [  85] = rx_phy_postflop_0 [  88];
  assign rx_upstream_data    [  86] = rx_phy_postflop_0 [  89];
  assign rx_upstream_data    [  87] = rx_phy_postflop_0 [  90];
  assign rx_upstream_data    [  88] = rx_phy_postflop_0 [  91];
  assign rx_upstream_data    [  89] = rx_phy_postflop_0 [  92];
  assign rx_upstream_data    [  90] = rx_phy_postflop_0 [  93];
  assign rx_upstream_data    [  91] = rx_phy_postflop_0 [  94];
  assign rx_upstream_data    [  92] = rx_phy_postflop_0 [  95];
  assign rx_upstream_data    [  93] = rx_phy_postflop_0 [  96];
  assign rx_upstream_data    [  94] = rx_phy_postflop_0 [  97];
  assign rx_upstream_data    [  95] = rx_phy_postflop_0 [  98];
  assign rx_upstream_data    [  96] = rx_phy_postflop_0 [  99];
  assign rx_upstream_data    [  97] = rx_phy_postflop_0 [ 100];
  assign rx_upstream_data    [  98] = rx_phy_postflop_0 [ 101];
  assign rx_upstream_data    [  99] = rx_phy_postflop_0 [ 102];
  assign rx_upstream_data    [ 100] = rx_phy_postflop_0 [ 103];
  assign rx_upstream_data    [ 101] = rx_phy_postflop_0 [ 104];
  assign rx_upstream_data    [ 102] = rx_phy_postflop_0 [ 105];
  assign rx_upstream_data    [ 103] = rx_phy_postflop_0 [ 106];
  assign rx_upstream_data    [ 104] = rx_phy_postflop_0 [ 107];
  assign rx_upstream_data    [ 105] = rx_phy_postflop_0 [ 108];
  assign rx_upstream_data    [ 106] = rx_phy_postflop_0 [ 109];
  assign rx_upstream_data    [ 107] = rx_phy_postflop_0 [ 110];
  assign rx_upstream_data    [ 108] = rx_phy_postflop_0 [ 111];
  assign rx_upstream_data    [ 109] = rx_phy_postflop_0 [ 112];
  assign rx_upstream_data    [ 110] = rx_phy_postflop_0 [ 113];
  assign rx_upstream_data    [ 111] = rx_phy_postflop_0 [ 114];
  assign rx_upstream_data    [ 112] = rx_phy_postflop_0 [ 115];
  assign rx_upstream_data    [ 113] = rx_phy_postflop_0 [ 116];
  assign rx_upstream_data    [ 114] = rx_phy_postflop_0 [ 117];
  assign rx_upstream_data    [ 115] = rx_phy_postflop_0 [ 118];
  assign rx_upstream_data    [ 116] = rx_phy_postflop_0 [ 119];
  assign rx_upstream_data    [ 117] = rx_phy_postflop_0 [ 120];
  assign rx_upstream_data    [ 118] = rx_phy_postflop_0 [ 121];
  assign rx_upstream_data    [ 119] = rx_phy_postflop_0 [ 122];
  assign rx_upstream_data    [ 120] = rx_phy_postflop_0 [ 123];
  assign rx_upstream_data    [ 121] = rx_phy_postflop_0 [ 124];
  assign rx_upstream_data    [ 122] = rx_phy_postflop_0 [ 125];
  assign rx_upstream_data    [ 123] = rx_phy_postflop_0 [ 126];
  assign rx_upstream_data    [ 124] = rx_phy_postflop_0 [ 127];
  assign rx_upstream_data    [ 125] = rx_phy_postflop_0 [ 128];
  assign rx_upstream_data    [ 126] = rx_phy_postflop_0 [ 129];
  assign rx_upstream_data    [ 127] = rx_phy_postflop_0 [ 130];
  assign rx_upstream_data    [ 128] = rx_phy_postflop_0 [ 131];
  assign rx_upstream_data    [ 129] = rx_phy_postflop_0 [ 132];
  assign rx_upstream_data    [ 130] = rx_phy_postflop_0 [ 133];
  assign rx_upstream_data    [ 131] = rx_phy_postflop_0 [ 134];
  assign rx_upstream_data    [ 132] = rx_phy_postflop_0 [ 135];
  assign rx_upstream_data    [ 133] = rx_phy_postflop_0 [ 136];
  assign rx_upstream_data    [ 134] = rx_phy_postflop_0 [ 137];
  assign rx_upstream_data    [ 135] = rx_phy_postflop_0 [ 138];
  assign rx_upstream_data    [ 136] = rx_phy_postflop_0 [ 139];
  assign rx_upstream_data    [ 137] = rx_phy_postflop_0 [ 140];
  assign rx_upstream_data    [ 138] = rx_phy_postflop_0 [ 141];
  assign rx_upstream_data    [ 139] = rx_phy_postflop_0 [ 142];
  assign rx_upstream_data    [ 140] = rx_phy_postflop_0 [ 143];
  assign rx_upstream_data    [ 141] = rx_phy_postflop_0 [ 144];
  assign rx_upstream_data    [ 142] = rx_phy_postflop_0 [ 145];
  assign rx_upstream_data    [ 143] = rx_phy_postflop_0 [ 146];
  assign rx_upstream_data    [ 144] = rx_phy_postflop_0 [ 147];
  assign rx_upstream_data    [ 145] = rx_phy_postflop_0 [ 148];
  assign rx_upstream_data    [ 146] = rx_phy_postflop_0 [ 149];
  assign rx_upstream_data    [ 147] = rx_phy_postflop_0 [ 150];
  assign rx_upstream_data    [ 148] = rx_phy_postflop_0 [ 151];
  assign rx_upstream_data    [ 149] = rx_phy_postflop_0 [ 152];
  assign rx_upstream_data    [ 150] = rx_phy_postflop_0 [ 153];
  assign rx_upstream_data    [ 151] = rx_phy_postflop_0 [ 154];
  assign rx_upstream_data    [ 152] = rx_phy_postflop_0 [ 155];
  assign rx_upstream_data    [ 153] = rx_phy_postflop_0 [ 156];
  assign rx_upstream_data    [ 154] = rx_phy_postflop_0 [ 157];
  assign rx_upstream_data    [ 155] = rx_phy_postflop_0 [ 158];
  assign rx_upstream_data    [ 156] = rx_phy_postflop_0 [ 159];
  assign rx_upstream_data    [ 157] = rx_phy_postflop_1 [   0];
  assign rx_upstream_data    [ 158] = rx_phy_postflop_1 [   1];
  assign rx_upstream_data    [ 159] = rx_phy_postflop_1 [   2];
  assign rx_upstream_data    [ 160] = rx_phy_postflop_1 [   3];
//       MARKER                     = rx_phy_postflop_1 [   4]
  assign rx_upstream_data    [ 161] = rx_phy_postflop_1 [   5];
  assign rx_upstream_data    [ 162] = rx_phy_postflop_1 [   6];
  assign rx_upstream_data    [ 163] = rx_phy_postflop_1 [   7];
  assign rx_upstream_data    [ 164] = rx_phy_postflop_1 [   8];
  assign rx_upstream_data    [ 165] = rx_phy_postflop_1 [   9];
  assign rx_upstream_data    [ 166] = rx_phy_postflop_1 [  10];
  assign rx_upstream_data    [ 167] = rx_phy_postflop_1 [  11];
  assign rx_upstream_data    [ 168] = rx_phy_postflop_1 [  12];
  assign rx_upstream_data    [ 169] = rx_phy_postflop_1 [  13];
  assign rx_upstream_data    [ 170] = rx_phy_postflop_1 [  14];
  assign rx_upstream_data    [ 171] = rx_phy_postflop_1 [  15];
  assign rx_upstream_data    [ 172] = rx_phy_postflop_1 [  16];
  assign rx_upstream_data    [ 173] = rx_phy_postflop_1 [  17];
  assign rx_upstream_data    [ 174] = rx_phy_postflop_1 [  18];
  assign rx_upstream_data    [ 175] = rx_phy_postflop_1 [  19];
  assign rx_upstream_data    [ 176] = rx_phy_postflop_1 [  20];
  assign rx_upstream_data    [ 177] = rx_phy_postflop_1 [  21];
  assign rx_upstream_data    [ 178] = rx_phy_postflop_1 [  22];
  assign rx_upstream_data    [ 179] = rx_phy_postflop_1 [  23];
  assign rx_upstream_data    [ 180] = rx_phy_postflop_1 [  24];
  assign rx_upstream_data    [ 181] = rx_phy_postflop_1 [  25];
  assign rx_upstream_data    [ 182] = rx_phy_postflop_1 [  26];
  assign rx_upstream_data    [ 183] = rx_phy_postflop_1 [  27];
  assign rx_upstream_data    [ 184] = rx_phy_postflop_1 [  28];
  assign rx_upstream_data    [ 185] = rx_phy_postflop_1 [  29];
  assign rx_upstream_data    [ 186] = rx_phy_postflop_1 [  30];
  assign rx_upstream_data    [ 187] = rx_phy_postflop_1 [  31];
  assign rx_upstream_data    [ 188] = rx_phy_postflop_1 [  32];
  assign rx_upstream_data    [ 189] = rx_phy_postflop_1 [  33];
  assign rx_upstream_data    [ 190] = rx_phy_postflop_1 [  34];
  assign rx_upstream_data    [ 191] = rx_phy_postflop_1 [  35];
  assign rx_upstream_data    [ 192] = rx_phy_postflop_1 [  36];
  assign rx_upstream_data    [ 193] = rx_phy_postflop_1 [  37];
  assign rx_upstream_data    [ 194] = rx_phy_postflop_1 [  38];
  assign rx_upstream_data    [ 195] = rx_phy_postflop_1 [  39];
  assign rx_upstream_data    [ 196] = rx_phy_postflop_1 [  40];
  assign rx_upstream_data    [ 197] = rx_phy_postflop_1 [  41];
  assign rx_upstream_data    [ 198] = rx_phy_postflop_1 [  42];
  assign rx_upstream_data    [ 199] = rx_phy_postflop_1 [  43];
  assign rx_upstream_data    [ 200] = rx_phy_postflop_1 [  44];
  assign rx_upstream_data    [ 201] = rx_phy_postflop_1 [  45];
  assign rx_upstream_data    [ 202] = rx_phy_postflop_1 [  46];
  assign rx_upstream_data    [ 203] = rx_phy_postflop_1 [  47];
  assign rx_upstream_data    [ 204] = rx_phy_postflop_1 [  48];
  assign rx_upstream_data    [ 205] = rx_phy_postflop_1 [  49];
  assign rx_upstream_data    [ 206] = rx_phy_postflop_1 [  50];
  assign rx_upstream_data    [ 207] = rx_phy_postflop_1 [  51];
  assign rx_upstream_data    [ 208] = rx_phy_postflop_1 [  52];
  assign rx_upstream_data    [ 209] = rx_phy_postflop_1 [  53];
  assign rx_upstream_data    [ 210] = rx_phy_postflop_1 [  54];
  assign rx_upstream_data    [ 211] = rx_phy_postflop_1 [  55];
  assign rx_upstream_data    [ 212] = rx_phy_postflop_1 [  56];
  assign rx_upstream_data    [ 213] = rx_phy_postflop_1 [  57];
  assign rx_upstream_data    [ 214] = rx_phy_postflop_1 [  58];
  assign rx_upstream_data    [ 215] = rx_phy_postflop_1 [  59];
  assign rx_upstream_data    [ 216] = rx_phy_postflop_1 [  60];
  assign rx_upstream_data    [ 217] = rx_phy_postflop_1 [  61];
  assign rx_upstream_data    [ 218] = rx_phy_postflop_1 [  62];
  assign rx_upstream_data    [ 219] = rx_phy_postflop_1 [  63];
  assign rx_upstream_data    [ 220] = rx_phy_postflop_1 [  64];
  assign rx_upstream_data    [ 221] = rx_phy_postflop_1 [  65];
  assign rx_upstream_data    [ 222] = rx_phy_postflop_1 [  66];
  assign rx_upstream_data    [ 223] = rx_phy_postflop_1 [  67];
  assign rx_upstream_data    [ 224] = rx_phy_postflop_1 [  68];
  assign rx_upstream_data    [ 225] = rx_phy_postflop_1 [  69];
  assign rx_upstream_data    [ 226] = rx_phy_postflop_1 [  70];
  assign rx_upstream_data    [ 227] = rx_phy_postflop_1 [  71];
  assign rx_upstream_data    [ 228] = rx_phy_postflop_1 [  72];
  assign rx_upstream_data    [ 229] = rx_phy_postflop_1 [  73];
  assign rx_upstream_data    [ 230] = rx_phy_postflop_1 [  74];
  assign rx_upstream_data    [ 231] = rx_phy_postflop_1 [  75];
//       STROBE                     = rx_phy_postflop_1 [  76]
  assign rx_upstream_data    [ 232] = rx_phy_postflop_1 [  77];
  assign rx_upstream_data    [ 233] = rx_phy_postflop_1 [  78];
  assign rx_upstream_data    [ 234] = rx_phy_postflop_1 [  79];
  assign rx_upstream_data    [ 235] = rx_phy_postflop_1 [  80];
  assign rx_upstream_data    [ 236] = rx_phy_postflop_1 [  81];
  assign rx_upstream_data    [ 237] = rx_phy_postflop_1 [  82];
  assign rx_upstream_data    [ 238] = rx_phy_postflop_1 [  83];
//       MARKER                     = rx_phy_postflop_1 [  84]
  assign rx_upstream_data    [ 239] = rx_phy_postflop_1 [  85];
  assign rx_upstream_data    [ 240] = rx_phy_postflop_1 [  86];
  assign rx_upstream_data    [ 241] = rx_phy_postflop_1 [  87];
  assign rx_upstream_data    [ 242] = rx_phy_postflop_1 [  88];
  assign rx_upstream_data    [ 243] = rx_phy_postflop_1 [  89];
  assign rx_upstream_data    [ 244] = rx_phy_postflop_1 [  90];
  assign rx_upstream_data    [ 245] = rx_phy_postflop_1 [  91];
  assign rx_upstream_data    [ 246] = rx_phy_postflop_1 [  92];
  assign rx_upstream_data    [ 247] = rx_phy_postflop_1 [  93];
  assign rx_upstream_data    [ 248] = rx_phy_postflop_1 [  94];
  assign rx_upstream_data    [ 249] = rx_phy_postflop_1 [  95];
  assign rx_upstream_data    [ 250] = rx_phy_postflop_1 [  96];
  assign rx_upstream_data    [ 251] = rx_phy_postflop_1 [  97];
  assign rx_upstream_data    [ 252] = rx_phy_postflop_1 [  98];
  assign rx_upstream_data    [ 253] = rx_phy_postflop_1 [  99];
  assign rx_upstream_data    [ 254] = rx_phy_postflop_1 [ 100];
  assign rx_upstream_data    [ 255] = rx_phy_postflop_1 [ 101];
  assign rx_upstream_data    [ 256] = rx_phy_postflop_1 [ 102];
  assign rx_upstream_data    [ 257] = rx_phy_postflop_1 [ 103];
  assign rx_upstream_data    [ 258] = rx_phy_postflop_1 [ 104];
  assign rx_upstream_data    [ 259] = rx_phy_postflop_1 [ 105];
  assign rx_upstream_data    [ 260] = rx_phy_postflop_1 [ 106];
  assign rx_upstream_data    [ 261] = rx_phy_postflop_1 [ 107];
  assign rx_upstream_data    [ 262] = rx_phy_postflop_1 [ 108];
  assign rx_upstream_data    [ 263] = rx_phy_postflop_1 [ 109];
  assign rx_upstream_data    [ 264] = rx_phy_postflop_1 [ 110];
  assign rx_upstream_data    [ 265] = rx_phy_postflop_1 [ 111];
  assign rx_upstream_data    [ 266] = rx_phy_postflop_1 [ 112];
  assign rx_upstream_data    [ 267] = rx_phy_postflop_1 [ 113];
  assign rx_upstream_data    [ 268] = rx_phy_postflop_1 [ 114];
  assign rx_upstream_data    [ 269] = rx_phy_postflop_1 [ 115];
  assign rx_upstream_data    [ 270] = rx_phy_postflop_1 [ 116];
  assign rx_upstream_data    [ 271] = rx_phy_postflop_1 [ 117];
  assign rx_upstream_data    [ 272] = rx_phy_postflop_1 [ 118];
  assign rx_upstream_data    [ 273] = rx_phy_postflop_1 [ 119];
  assign rx_upstream_data    [ 274] = rx_phy_postflop_1 [ 120];
  assign rx_upstream_data    [ 275] = rx_phy_postflop_1 [ 121];
  assign rx_upstream_data    [ 276] = rx_phy_postflop_1 [ 122];
  assign rx_upstream_data    [ 277] = rx_phy_postflop_1 [ 123];
  assign rx_upstream_data    [ 278] = rx_phy_postflop_1 [ 124];
  assign rx_upstream_data    [ 279] = rx_phy_postflop_1 [ 125];
  assign rx_upstream_data    [ 280] = rx_phy_postflop_1 [ 126];
  assign rx_upstream_data    [ 281] = rx_phy_postflop_1 [ 127];
  assign rx_upstream_data    [ 282] = rx_phy_postflop_1 [ 128];
  assign rx_upstream_data    [ 283] = rx_phy_postflop_1 [ 129];
  assign rx_upstream_data    [ 284] = rx_phy_postflop_1 [ 130];
  assign rx_upstream_data    [ 285] = rx_phy_postflop_1 [ 131];
  assign rx_upstream_data    [ 286] = rx_phy_postflop_1 [ 132];
  assign rx_upstream_data    [ 287] = rx_phy_postflop_1 [ 133];
  assign rx_upstream_data    [ 288] = rx_phy_postflop_1 [ 134];
  assign rx_upstream_data    [ 289] = rx_phy_postflop_1 [ 135];
  assign rx_upstream_data    [ 290] = rx_phy_postflop_1 [ 136];
  assign rx_upstream_data    [ 291] = rx_phy_postflop_1 [ 137];
  assign rx_upstream_data    [ 292] = rx_phy_postflop_1 [ 138];
  assign rx_upstream_data    [ 293] = rx_phy_postflop_1 [ 139];
  assign rx_upstream_data    [ 294] = rx_phy_postflop_1 [ 140];
  assign rx_upstream_data    [ 295] = rx_phy_postflop_1 [ 141];
  assign rx_upstream_data    [ 296] = rx_phy_postflop_1 [ 142];
  assign rx_upstream_data    [ 297] = rx_phy_postflop_1 [ 143];
  assign rx_upstream_data    [ 298] = rx_phy_postflop_1 [ 144];
  assign rx_upstream_data    [ 299] = rx_phy_postflop_1 [ 145];
  assign rx_upstream_data    [ 300] = rx_phy_postflop_1 [ 146];
  assign rx_upstream_data    [ 301] = rx_phy_postflop_1 [ 147];
  assign rx_upstream_data    [ 302] = rx_phy_postflop_1 [ 148];
  assign rx_upstream_data    [ 303] = rx_phy_postflop_1 [ 149];
  assign rx_upstream_data    [ 304] = rx_phy_postflop_1 [ 150];
  assign rx_upstream_data    [ 305] = rx_phy_postflop_1 [ 151];
  assign rx_upstream_data    [ 306] = rx_phy_postflop_1 [ 152];
  assign rx_upstream_data    [ 307] = rx_phy_postflop_1 [ 153];
  assign rx_upstream_data    [ 308] = rx_phy_postflop_1 [ 154];
  assign rx_upstream_data    [ 309] = rx_phy_postflop_1 [ 155];
  assign rx_upstream_data    [ 310] = rx_phy_postflop_1 [ 156];
  assign rx_upstream_data    [ 311] = rx_phy_postflop_1 [ 157];
  assign rx_upstream_data    [ 312] = rx_phy_postflop_1 [ 158];
  assign rx_upstream_data    [ 313] = rx_phy_postflop_1 [ 159];
  assign rx_upstream_data    [ 314] = rx_phy_postflop_2 [   0];
  assign rx_upstream_data    [ 315] = rx_phy_postflop_2 [   1];
  assign rx_upstream_data    [ 316] = rx_phy_postflop_2 [   2];
  assign rx_upstream_data    [ 317] = rx_phy_postflop_2 [   3];
//       MARKER                     = rx_phy_postflop_2 [   4]
  assign rx_upstream_data    [ 318] = rx_phy_postflop_2 [   5];
  assign rx_upstream_data    [ 319] = rx_phy_postflop_2 [   6];
  assign rx_upstream_data    [ 320] = rx_phy_postflop_2 [   7];
  assign rx_upstream_data    [ 321] = rx_phy_postflop_2 [   8];
  assign rx_upstream_data    [ 322] = rx_phy_postflop_2 [   9];
  assign rx_upstream_data    [ 323] = rx_phy_postflop_2 [  10];
  assign rx_upstream_data    [ 324] = rx_phy_postflop_2 [  11];
  assign rx_upstream_data    [ 325] = rx_phy_postflop_2 [  12];
  assign rx_upstream_data    [ 326] = rx_phy_postflop_2 [  13];
  assign rx_upstream_data    [ 327] = rx_phy_postflop_2 [  14];
  assign rx_upstream_data    [ 328] = rx_phy_postflop_2 [  15];
  assign rx_upstream_data    [ 329] = rx_phy_postflop_2 [  16];
  assign rx_upstream_data    [ 330] = rx_phy_postflop_2 [  17];
  assign rx_upstream_data    [ 331] = rx_phy_postflop_2 [  18];
  assign rx_upstream_data    [ 332] = rx_phy_postflop_2 [  19];
  assign rx_upstream_data    [ 333] = rx_phy_postflop_2 [  20];
  assign rx_upstream_data    [ 334] = rx_phy_postflop_2 [  21];
  assign rx_upstream_data    [ 335] = rx_phy_postflop_2 [  22];
  assign rx_upstream_data    [ 336] = rx_phy_postflop_2 [  23];
  assign rx_upstream_data    [ 337] = rx_phy_postflop_2 [  24];
  assign rx_upstream_data    [ 338] = rx_phy_postflop_2 [  25];
  assign rx_upstream_data    [ 339] = rx_phy_postflop_2 [  26];
  assign rx_upstream_data    [ 340] = rx_phy_postflop_2 [  27];
  assign rx_upstream_data    [ 341] = rx_phy_postflop_2 [  28];
  assign rx_upstream_data    [ 342] = rx_phy_postflop_2 [  29];
  assign rx_upstream_data    [ 343] = rx_phy_postflop_2 [  30];
  assign rx_upstream_data    [ 344] = rx_phy_postflop_2 [  31];
  assign rx_upstream_data    [ 345] = rx_phy_postflop_2 [  32];
  assign rx_upstream_data    [ 346] = rx_phy_postflop_2 [  33];
  assign rx_upstream_data    [ 347] = rx_phy_postflop_2 [  34];
  assign rx_upstream_data    [ 348] = rx_phy_postflop_2 [  35];
  assign rx_upstream_data    [ 349] = rx_phy_postflop_2 [  36];
  assign rx_upstream_data    [ 350] = rx_phy_postflop_2 [  37];
  assign rx_upstream_data    [ 351] = rx_phy_postflop_2 [  38];
  assign rx_upstream_data    [ 352] = rx_phy_postflop_2 [  39];
  assign rx_upstream_data    [ 353] = rx_phy_postflop_2 [  40];
  assign rx_upstream_data    [ 354] = rx_phy_postflop_2 [  41];
  assign rx_upstream_data    [ 355] = rx_phy_postflop_2 [  42];
  assign rx_upstream_data    [ 356] = rx_phy_postflop_2 [  43];
  assign rx_upstream_data    [ 357] = rx_phy_postflop_2 [  44];
  assign rx_upstream_data    [ 358] = rx_phy_postflop_2 [  45];
  assign rx_upstream_data    [ 359] = rx_phy_postflop_2 [  46];
  assign rx_upstream_data    [ 360] = rx_phy_postflop_2 [  47];
  assign rx_upstream_data    [ 361] = rx_phy_postflop_2 [  48];
  assign rx_upstream_data    [ 362] = rx_phy_postflop_2 [  49];
  assign rx_upstream_data    [ 363] = rx_phy_postflop_2 [  50];
  assign rx_upstream_data    [ 364] = rx_phy_postflop_2 [  51];
  assign rx_upstream_data    [ 365] = rx_phy_postflop_2 [  52];
  assign rx_upstream_data    [ 366] = rx_phy_postflop_2 [  53];
  assign rx_upstream_data    [ 367] = rx_phy_postflop_2 [  54];
  assign rx_upstream_data    [ 368] = rx_phy_postflop_2 [  55];
  assign rx_upstream_data    [ 369] = rx_phy_postflop_2 [  56];
  assign rx_upstream_data    [ 370] = rx_phy_postflop_2 [  57];
  assign rx_upstream_data    [ 371] = rx_phy_postflop_2 [  58];
  assign rx_upstream_data    [ 372] = rx_phy_postflop_2 [  59];
  assign rx_upstream_data    [ 373] = rx_phy_postflop_2 [  60];
  assign rx_upstream_data    [ 374] = rx_phy_postflop_2 [  61];
  assign rx_upstream_data    [ 375] = rx_phy_postflop_2 [  62];
  assign rx_upstream_data    [ 376] = rx_phy_postflop_2 [  63];
  assign rx_upstream_data    [ 377] = rx_phy_postflop_2 [  64];
  assign rx_upstream_data    [ 378] = rx_phy_postflop_2 [  65];
  assign rx_upstream_data    [ 379] = rx_phy_postflop_2 [  66];
  assign rx_upstream_data    [ 380] = rx_phy_postflop_2 [  67];
  assign rx_upstream_data    [ 381] = rx_phy_postflop_2 [  68];
  assign rx_upstream_data    [ 382] = rx_phy_postflop_2 [  69];
  assign rx_upstream_data    [ 383] = rx_phy_postflop_2 [  70];
  assign rx_upstream_data    [ 384] = rx_phy_postflop_2 [  71];
  assign rx_upstream_data    [ 385] = rx_phy_postflop_2 [  72];
  assign rx_upstream_data    [ 386] = rx_phy_postflop_2 [  73];
  assign rx_upstream_data    [ 387] = rx_phy_postflop_2 [  74];
  assign rx_upstream_data    [ 388] = rx_phy_postflop_2 [  75];
//       STROBE                     = rx_phy_postflop_2 [  76]
  assign rx_upstream_data    [ 389] = rx_phy_postflop_2 [  77];
  assign rx_upstream_data    [ 390] = rx_phy_postflop_2 [  78];
  assign rx_upstream_data    [ 391] = rx_phy_postflop_2 [  79];
  assign rx_upstream_data    [ 392] = rx_phy_postflop_2 [  80];
  assign rx_upstream_data    [ 393] = rx_phy_postflop_2 [  81];
  assign rx_upstream_data    [ 394] = rx_phy_postflop_2 [  82];
  assign rx_upstream_data    [ 395] = rx_phy_postflop_2 [  83];
//       MARKER                     = rx_phy_postflop_2 [  84]
  assign rx_upstream_data    [ 396] = rx_phy_postflop_2 [  85];
  assign rx_upstream_data    [ 397] = rx_phy_postflop_2 [  86];
  assign rx_upstream_data    [ 398] = rx_phy_postflop_2 [  87];
  assign rx_upstream_data    [ 399] = rx_phy_postflop_2 [  88];
  assign rx_upstream_data    [ 400] = rx_phy_postflop_2 [  89];
  assign rx_upstream_data    [ 401] = rx_phy_postflop_2 [  90];
  assign rx_upstream_data    [ 402] = rx_phy_postflop_2 [  91];
  assign rx_upstream_data    [ 403] = rx_phy_postflop_2 [  92];
  assign rx_upstream_data    [ 404] = rx_phy_postflop_2 [  93];
  assign rx_upstream_data    [ 405] = rx_phy_postflop_2 [  94];
  assign rx_upstream_data    [ 406] = rx_phy_postflop_2 [  95];
  assign rx_upstream_data    [ 407] = rx_phy_postflop_2 [  96];
  assign rx_upstream_data    [ 408] = rx_phy_postflop_2 [  97];
  assign rx_upstream_data    [ 409] = rx_phy_postflop_2 [  98];
  assign rx_upstream_data    [ 410] = rx_phy_postflop_2 [  99];
  assign rx_upstream_data    [ 411] = rx_phy_postflop_2 [ 100];
  assign rx_upstream_data    [ 412] = rx_phy_postflop_2 [ 101];
  assign rx_upstream_data    [ 413] = rx_phy_postflop_2 [ 102];
  assign rx_upstream_data    [ 414] = rx_phy_postflop_2 [ 103];
  assign rx_upstream_data    [ 415] = rx_phy_postflop_2 [ 104];
  assign rx_upstream_data    [ 416] = rx_phy_postflop_2 [ 105];
  assign rx_upstream_data    [ 417] = rx_phy_postflop_2 [ 106];
  assign rx_upstream_data    [ 418] = rx_phy_postflop_2 [ 107];
  assign rx_upstream_data    [ 419] = rx_phy_postflop_2 [ 108];
  assign rx_upstream_data    [ 420] = rx_phy_postflop_2 [ 109];
  assign rx_upstream_data    [ 421] = rx_phy_postflop_2 [ 110];
  assign rx_upstream_data    [ 422] = rx_phy_postflop_2 [ 111];
  assign rx_upstream_data    [ 423] = rx_phy_postflop_2 [ 112];
  assign rx_upstream_data    [ 424] = rx_phy_postflop_2 [ 113];
  assign rx_upstream_data    [ 425] = rx_phy_postflop_2 [ 114];
  assign rx_upstream_data    [ 426] = rx_phy_postflop_2 [ 115];
  assign rx_upstream_data    [ 427] = rx_phy_postflop_2 [ 116];
  assign rx_upstream_data    [ 428] = rx_phy_postflop_2 [ 117];
  assign rx_upstream_data    [ 429] = rx_phy_postflop_2 [ 118];
  assign rx_upstream_data    [ 430] = rx_phy_postflop_2 [ 119];
  assign rx_upstream_data    [ 431] = rx_phy_postflop_2 [ 120];
  assign rx_upstream_data    [ 432] = rx_phy_postflop_2 [ 121];
  assign rx_upstream_data    [ 433] = rx_phy_postflop_2 [ 122];
  assign rx_upstream_data    [ 434] = rx_phy_postflop_2 [ 123];
  assign rx_upstream_data    [ 435] = rx_phy_postflop_2 [ 124];
  assign rx_upstream_data    [ 436] = rx_phy_postflop_2 [ 125];
  assign rx_upstream_data    [ 437] = rx_phy_postflop_2 [ 126];
  assign rx_upstream_data    [ 438] = rx_phy_postflop_2 [ 127];
  assign rx_upstream_data    [ 439] = rx_phy_postflop_2 [ 128];
  assign rx_upstream_data    [ 440] = rx_phy_postflop_2 [ 129];
  assign rx_upstream_data    [ 441] = rx_phy_postflop_2 [ 130];
  assign rx_upstream_data    [ 442] = rx_phy_postflop_2 [ 131];
  assign rx_upstream_data    [ 443] = rx_phy_postflop_2 [ 132];
  assign rx_upstream_data    [ 444] = rx_phy_postflop_2 [ 133];
  assign rx_upstream_data    [ 445] = rx_phy_postflop_2 [ 134];
  assign rx_upstream_data    [ 446] = rx_phy_postflop_2 [ 135];
  assign rx_upstream_data    [ 447] = rx_phy_postflop_2 [ 136];
  assign rx_upstream_data    [ 448] = rx_phy_postflop_2 [ 137];
  assign rx_upstream_data    [ 449] = rx_phy_postflop_2 [ 138];
  assign rx_upstream_data    [ 450] = rx_phy_postflop_2 [ 139];
  assign rx_upstream_data    [ 451] = rx_phy_postflop_2 [ 140];
  assign rx_upstream_data    [ 452] = rx_phy_postflop_2 [ 141];
  assign rx_upstream_data    [ 453] = rx_phy_postflop_2 [ 142];
  assign rx_upstream_data    [ 454] = rx_phy_postflop_2 [ 143];
  assign rx_upstream_data    [ 455] = rx_phy_postflop_2 [ 144];
  assign rx_upstream_data    [ 456] = rx_phy_postflop_2 [ 145];
  assign rx_upstream_data    [ 457] = rx_phy_postflop_2 [ 146];
  assign rx_upstream_data    [ 458] = rx_phy_postflop_2 [ 147];
  assign rx_upstream_data    [ 459] = rx_phy_postflop_2 [ 148];
  assign rx_upstream_data    [ 460] = rx_phy_postflop_2 [ 149];
  assign rx_upstream_data    [ 461] = rx_phy_postflop_2 [ 150];
  assign rx_upstream_data    [ 462] = rx_phy_postflop_2 [ 151];
  assign rx_upstream_data    [ 463] = rx_phy_postflop_2 [ 152];
  assign rx_upstream_data    [ 464] = rx_phy_postflop_2 [ 153];
  assign rx_upstream_data    [ 465] = rx_phy_postflop_2 [ 154];
  assign rx_upstream_data    [ 466] = rx_phy_postflop_2 [ 155];
  assign rx_upstream_data    [ 467] = rx_phy_postflop_2 [ 156];
  assign rx_upstream_data    [ 468] = rx_phy_postflop_2 [ 157];
  assign rx_upstream_data    [ 469] = rx_phy_postflop_2 [ 158];
  assign rx_upstream_data    [ 470] = rx_phy_postflop_2 [ 159];
  assign rx_upstream_data    [ 471] = rx_phy_postflop_3 [   0];
  assign rx_upstream_data    [ 472] = rx_phy_postflop_3 [   1];
  assign rx_upstream_data    [ 473] = rx_phy_postflop_3 [   2];
  assign rx_upstream_data    [ 474] = rx_phy_postflop_3 [   3];
//       MARKER                     = rx_phy_postflop_3 [   4]
  assign rx_upstream_data    [ 475] = rx_phy_postflop_3 [   5];
  assign rx_upstream_data    [ 476] = rx_phy_postflop_3 [   6];
  assign rx_upstream_data    [ 477] = rx_phy_postflop_3 [   7];
  assign rx_upstream_data    [ 478] = rx_phy_postflop_3 [   8];
  assign rx_upstream_data    [ 479] = rx_phy_postflop_3 [   9];
  assign rx_upstream_data    [ 480] = rx_phy_postflop_3 [  10];
  assign rx_upstream_data    [ 481] = rx_phy_postflop_3 [  11];
  assign rx_upstream_data    [ 482] = rx_phy_postflop_3 [  12];
  assign rx_upstream_data    [ 483] = rx_phy_postflop_3 [  13];
  assign rx_upstream_data    [ 484] = rx_phy_postflop_3 [  14];
  assign rx_upstream_data    [ 485] = rx_phy_postflop_3 [  15];
  assign rx_upstream_data    [ 486] = rx_phy_postflop_3 [  16];
  assign rx_upstream_data    [ 487] = rx_phy_postflop_3 [  17];
  assign rx_upstream_data    [ 488] = rx_phy_postflop_3 [  18];
  assign rx_upstream_data    [ 489] = rx_phy_postflop_3 [  19];
  assign rx_upstream_data    [ 490] = rx_phy_postflop_3 [  20];
  assign rx_upstream_data    [ 491] = rx_phy_postflop_3 [  21];
  assign rx_upstream_data    [ 492] = rx_phy_postflop_3 [  22];
  assign rx_upstream_data    [ 493] = rx_phy_postflop_3 [  23];
  assign rx_upstream_data    [ 494] = rx_phy_postflop_3 [  24];
  assign rx_upstream_data    [ 495] = rx_phy_postflop_3 [  25];
  assign rx_upstream_data    [ 496] = rx_phy_postflop_3 [  26];
  assign rx_upstream_data    [ 497] = rx_phy_postflop_3 [  27];
  assign rx_upstream_data    [ 498] = rx_phy_postflop_3 [  28];
  assign rx_upstream_data    [ 499] = rx_phy_postflop_3 [  29];
  assign rx_upstream_data    [ 500] = rx_phy_postflop_3 [  30];
  assign rx_upstream_data    [ 501] = rx_phy_postflop_3 [  31];
  assign rx_upstream_data    [ 502] = rx_phy_postflop_3 [  32];
  assign rx_upstream_data    [ 503] = rx_phy_postflop_3 [  33];
  assign rx_upstream_data    [ 504] = rx_phy_postflop_3 [  34];
  assign rx_upstream_data    [ 505] = rx_phy_postflop_3 [  35];
  assign rx_upstream_data    [ 506] = rx_phy_postflop_3 [  36];
  assign rx_upstream_data    [ 507] = rx_phy_postflop_3 [  37];
  assign rx_upstream_data    [ 508] = rx_phy_postflop_3 [  38];
  assign rx_upstream_data    [ 509] = rx_phy_postflop_3 [  39];
  assign rx_upstream_data    [ 510] = rx_phy_postflop_3 [  40];
  assign rx_upstream_data    [ 511] = rx_phy_postflop_3 [  41];
  assign rx_upstream_data    [ 512] = rx_phy_postflop_3 [  42];
  assign rx_upstream_data    [ 513] = rx_phy_postflop_3 [  43];
  assign rx_upstream_data    [ 514] = rx_phy_postflop_3 [  44];
  assign rx_upstream_data    [ 515] = rx_phy_postflop_3 [  45];
  assign rx_upstream_data    [ 516] = rx_phy_postflop_3 [  46];
  assign rx_upstream_data    [ 517] = rx_phy_postflop_3 [  47];
  assign rx_upstream_data    [ 518] = rx_phy_postflop_3 [  48];
  assign rx_upstream_data    [ 519] = rx_phy_postflop_3 [  49];
  assign rx_upstream_data    [ 520] = rx_phy_postflop_3 [  50];
  assign rx_upstream_data    [ 521] = rx_phy_postflop_3 [  51];
  assign rx_upstream_data    [ 522] = rx_phy_postflop_3 [  52];
  assign rx_upstream_data    [ 523] = rx_phy_postflop_3 [  53];
  assign rx_upstream_data    [ 524] = rx_phy_postflop_3 [  54];
  assign rx_upstream_data    [ 525] = rx_phy_postflop_3 [  55];
  assign rx_upstream_data    [ 526] = rx_phy_postflop_3 [  56];
  assign rx_upstream_data    [ 527] = rx_phy_postflop_3 [  57];
  assign rx_upstream_data    [ 528] = rx_phy_postflop_3 [  58];
  assign rx_upstream_data    [ 529] = rx_phy_postflop_3 [  59];
  assign rx_upstream_data    [ 530] = rx_phy_postflop_3 [  60];
  assign rx_upstream_data    [ 531] = rx_phy_postflop_3 [  61];
  assign rx_upstream_data    [ 532] = rx_phy_postflop_3 [  62];
  assign rx_upstream_data    [ 533] = rx_phy_postflop_3 [  63];
  assign rx_upstream_data    [ 534] = rx_phy_postflop_3 [  64];
  assign rx_upstream_data    [ 535] = rx_phy_postflop_3 [  65];
  assign rx_upstream_data    [ 536] = rx_phy_postflop_3 [  66];
  assign rx_upstream_data    [ 537] = rx_phy_postflop_3 [  67];
  assign rx_upstream_data    [ 538] = rx_phy_postflop_3 [  68];
  assign rx_upstream_data    [ 539] = rx_phy_postflop_3 [  69];
  assign rx_upstream_data    [ 540] = rx_phy_postflop_3 [  70];
  assign rx_upstream_data    [ 541] = rx_phy_postflop_3 [  71];
  assign rx_upstream_data    [ 542] = rx_phy_postflop_3 [  72];
  assign rx_upstream_data    [ 543] = rx_phy_postflop_3 [  73];
  assign rx_upstream_data    [ 544] = rx_phy_postflop_3 [  74];
  assign rx_upstream_data    [ 545] = rx_phy_postflop_3 [  75];
//       STROBE                     = rx_phy_postflop_3 [  76]
  assign rx_upstream_data    [ 546] = rx_phy_postflop_3 [  77];
  assign rx_upstream_data    [ 547] = rx_phy_postflop_3 [  78];
  assign rx_upstream_data    [ 548] = rx_phy_postflop_3 [  79];
  assign rx_upstream_data    [ 549] = rx_phy_postflop_3 [  80];
  assign rx_upstream_data    [ 550] = rx_phy_postflop_3 [  81];
  assign rx_upstream_data    [ 551] = rx_phy_postflop_3 [  82];
  assign rx_upstream_data    [ 552] = rx_phy_postflop_3 [  83];
//       MARKER                     = rx_phy_postflop_3 [  84]
  assign rx_upstream_data    [ 553] = rx_phy_postflop_3 [  85];
  assign rx_upstream_data    [ 554] = rx_phy_postflop_3 [  86];
  assign rx_upstream_data    [ 555] = rx_phy_postflop_3 [  87];
  assign rx_upstream_data    [ 556] = rx_phy_postflop_3 [  88];
  assign rx_upstream_data    [ 557] = rx_phy_postflop_3 [  89];
  assign rx_upstream_data    [ 558] = rx_phy_postflop_3 [  90];
  assign rx_upstream_data    [ 559] = rx_phy_postflop_3 [  91];
  assign rx_upstream_data    [ 560] = rx_phy_postflop_3 [  92];
  assign rx_upstream_data    [ 561] = rx_phy_postflop_3 [  93];
  assign rx_upstream_data    [ 562] = rx_phy_postflop_3 [  94];
  assign rx_upstream_data    [ 563] = rx_phy_postflop_3 [  95];
  assign rx_upstream_data    [ 564] = rx_phy_postflop_3 [  96];
  assign rx_upstream_data    [ 565] = rx_phy_postflop_3 [  97];
  assign rx_upstream_data    [ 566] = rx_phy_postflop_3 [  98];
  assign rx_upstream_data    [ 567] = rx_phy_postflop_3 [  99];
  assign rx_upstream_data    [ 568] = rx_phy_postflop_3 [ 100];
  assign rx_upstream_data    [ 569] = rx_phy_postflop_3 [ 101];
  assign rx_upstream_data    [ 570] = rx_phy_postflop_3 [ 102];
  assign rx_upstream_data    [ 571] = rx_phy_postflop_3 [ 103];
  assign rx_upstream_data    [ 572] = rx_phy_postflop_3 [ 104];
  assign rx_upstream_data    [ 573] = rx_phy_postflop_3 [ 105];
  assign rx_upstream_data    [ 574] = rx_phy_postflop_3 [ 106];
  assign rx_upstream_data    [ 575] = rx_phy_postflop_3 [ 107];
  assign rx_upstream_data    [ 576] = rx_phy_postflop_3 [ 108];
  assign rx_upstream_data    [ 577] = rx_phy_postflop_3 [ 109];
  assign rx_upstream_data    [ 578] = rx_phy_postflop_3 [ 110];
  assign rx_upstream_data    [ 579] = rx_phy_postflop_3 [ 111];
  assign rx_upstream_data    [ 580] = rx_phy_postflop_3 [ 112];
  assign rx_upstream_data    [ 581] = rx_phy_postflop_3 [ 113];
  assign rx_upstream_data    [ 582] = rx_phy_postflop_3 [ 114];
  assign rx_upstream_data    [ 583] = rx_phy_postflop_3 [ 115];
  assign rx_upstream_data    [ 584] = rx_phy_postflop_3 [ 116];
  assign rx_upstream_data    [ 585] = rx_phy_postflop_3 [ 117];
  assign rx_upstream_data    [ 586] = rx_phy_postflop_3 [ 118];
  assign rx_upstream_data    [ 587] = rx_phy_postflop_3 [ 119];
  assign rx_upstream_data    [ 588] = rx_phy_postflop_3 [ 120];
//       nc                         = rx_phy_postflop_3 [ 121];
//       nc                         = rx_phy_postflop_3 [ 122];
//       nc                         = rx_phy_postflop_3 [ 123];
//       nc                         = rx_phy_postflop_3 [ 124];
//       nc                         = rx_phy_postflop_3 [ 125];
//       nc                         = rx_phy_postflop_3 [ 126];
//       nc                         = rx_phy_postflop_3 [ 127];
//       nc                         = rx_phy_postflop_3 [ 128];
//       nc                         = rx_phy_postflop_3 [ 129];
//       nc                         = rx_phy_postflop_3 [ 130];
//       nc                         = rx_phy_postflop_3 [ 131];
//       nc                         = rx_phy_postflop_3 [ 132];
//       nc                         = rx_phy_postflop_3 [ 133];
//       nc                         = rx_phy_postflop_3 [ 134];
//       nc                         = rx_phy_postflop_3 [ 135];
//       nc                         = rx_phy_postflop_3 [ 136];
//       nc                         = rx_phy_postflop_3 [ 137];
//       nc                         = rx_phy_postflop_3 [ 138];
//       nc                         = rx_phy_postflop_3 [ 139];
//       nc                         = rx_phy_postflop_3 [ 140];
//       nc                         = rx_phy_postflop_3 [ 141];
//       nc                         = rx_phy_postflop_3 [ 142];
//       nc                         = rx_phy_postflop_3 [ 143];
//       nc                         = rx_phy_postflop_3 [ 144];
//       nc                         = rx_phy_postflop_3 [ 145];
//       nc                         = rx_phy_postflop_3 [ 146];
//       nc                         = rx_phy_postflop_3 [ 147];
//       nc                         = rx_phy_postflop_3 [ 148];
//       nc                         = rx_phy_postflop_3 [ 149];
//       nc                         = rx_phy_postflop_3 [ 150];
//       nc                         = rx_phy_postflop_3 [ 151];
//       nc                         = rx_phy_postflop_3 [ 152];
//       nc                         = rx_phy_postflop_3 [ 153];
//       nc                         = rx_phy_postflop_3 [ 154];
//       nc                         = rx_phy_postflop_3 [ 155];
//       nc                         = rx_phy_postflop_3 [ 156];
//       nc                         = rx_phy_postflop_3 [ 157];
//       nc                         = rx_phy_postflop_3 [ 158];
//       nc                         = rx_phy_postflop_3 [ 159];

// RX Section
//////////////////////////////////////////////////////////////////


endmodule
