`ifndef _CA_COVERAGE_
`define _CA_COVERAGE_
//////////////////////////////////////////////////////////////////

covergroup  ca_cfg_covergroup with function sample(ca_cfg_c  ca_cfg);

endgroup : ca_cfg_covergroup
    
//////////////////////////////////////////////////////////////////
`endif
