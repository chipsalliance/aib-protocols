////////////////////////////////////////////////////////////
//
//        (C) Copyright 2021 Eximius Design
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
////////////////////////////////////////////////////////////

module axi_st_d128_asym_quarter_slave_concat  (

// Data from Logic Links
  output logic [ 583:   0]   rx_st_data          ,
  output logic               rx_st_push_ovrd     ,
  output logic               rx_st_pushbit       ,
  input  logic [   3:   0]   tx_st_credit        ,

// PHY Interconnect
  output logic [ 319:   0]   tx_phy0             ,
  input  logic [ 319:   0]   rx_phy0             ,
  output logic [ 319:   0]   tx_phy1             ,
  input  logic [ 319:   0]   rx_phy1             ,

  input  logic               clk_wr              ,
  input  logic               clk_rd              ,
  input  logic               rst_wr_n            ,
  input  logic               rst_rd_n            ,

  input  logic               m_gen2_mode         ,
  input  logic               tx_online           ,

  input  logic               tx_stb_userbit      ,
  input  logic [   3:   0]   tx_mrk_userbit      

);

// No TX Packetization, so tie off packetization signals

// No RX Packetization, so tie off packetization signals
  assign rx_st_push_ovrd                    = 1'b0                               ;

//////////////////////////////////////////////////////////////////
// TX Section

//   TX_CH_WIDTH           = 320; // Gen2Only running at Quarter Rate
//   TX_DATA_WIDTH         = 296; // Usable Data per Channel
//   TX_PERSISTENT_STROBE  = 1'b1;
//   TX_PERSISTENT_MARKER  = 1'b1;
//   TX_STROBE_GEN2_LOC    = 'd1;
//   TX_MARKER_GEN2_LOC    = 'd0;
//   TX_STROBE_GEN1_LOC    = 'd38;
//   TX_MARKER_GEN1_LOC    = 'd39;
//   TX_ENABLE_STROBE      = 1'b1;
//   TX_ENABLE_MARKER      = 1'b1;
//   TX_DBI_PRESENT        = 1'b1;
//   TX_REG_PHY            = 1'b0;

  localparam TX_REG_PHY    = 1'b0;  // If set, this enables boundary FF for timing reasons

  logic [ 319:   0]                              tx_phy_preflop_0              ;
  logic [ 319:   0]                              tx_phy_preflop_1              ;
  logic [ 319:   0]                              tx_phy_flop_0_reg             ;
  logic [ 319:   0]                              tx_phy_flop_1_reg             ;

  always_ff @(posedge clk_wr or negedge rst_wr_n)
  if (~rst_wr_n)
  begin
    tx_phy_flop_0_reg                       <= 320'b0                                  ;
    tx_phy_flop_1_reg                       <= 320'b0                                  ;
  end
  else
  begin
    tx_phy_flop_0_reg                       <= tx_phy_preflop_0                        ;
    tx_phy_flop_1_reg                       <= tx_phy_preflop_1                        ;
  end

  assign tx_phy0                            = TX_REG_PHY ? tx_phy_flop_0_reg : tx_phy_preflop_0               ;
  assign tx_phy1                            = TX_REG_PHY ? tx_phy_flop_1_reg : tx_phy_preflop_1               ;

  logic                                          tx_st_credit_r0               ;
  logic                                          tx_st_credit_r1               ;
  logic                                          tx_st_credit_r2               ;
  logic                                          tx_st_credit_r3               ;

  // Asymmetric Credit Logic
  assign tx_st_credit_r0                    = tx_st_credit         [   0 +:   1] ;
  assign tx_st_credit_r1                    = tx_st_credit         [   1 +:   1] ;
  assign tx_st_credit_r2                    = tx_st_credit         [   2 +:   1] ;
  assign tx_st_credit_r3                    = tx_st_credit         [   3 +:   1] ;

  assign tx_phy_preflop_0 [   0] = tx_mrk_userbit[0]          ; // MARKER
  assign tx_phy_preflop_0 [   1] = tx_stb_userbit             ; // STROBE
  assign tx_phy_preflop_0 [   2] = tx_st_credit_r0            ;
  assign tx_phy_preflop_0 [   3] = 1'b0                       ;
  assign tx_phy_preflop_0 [   4] = 1'b0                       ;
  assign tx_phy_preflop_0 [   5] = 1'b0                       ;
  assign tx_phy_preflop_0 [   6] = 1'b0                       ;
  assign tx_phy_preflop_0 [   7] = 1'b0                       ;
  assign tx_phy_preflop_0 [   8] = 1'b0                       ;
  assign tx_phy_preflop_0 [   9] = 1'b0                       ;
  assign tx_phy_preflop_0 [  10] = 1'b0                       ;
  assign tx_phy_preflop_0 [  11] = 1'b0                       ;
  assign tx_phy_preflop_0 [  12] = 1'b0                       ;
  assign tx_phy_preflop_0 [  13] = 1'b0                       ;
  assign tx_phy_preflop_0 [  14] = 1'b0                       ;
  assign tx_phy_preflop_0 [  15] = 1'b0                       ;
  assign tx_phy_preflop_0 [  16] = 1'b0                       ;
  assign tx_phy_preflop_0 [  17] = 1'b0                       ;
  assign tx_phy_preflop_0 [  18] = 1'b0                       ;
  assign tx_phy_preflop_0 [  19] = 1'b0                       ;
  assign tx_phy_preflop_0 [  20] = 1'b0                       ;
  assign tx_phy_preflop_0 [  21] = 1'b0                       ;
  assign tx_phy_preflop_0 [  22] = 1'b0                       ;
  assign tx_phy_preflop_0 [  23] = 1'b0                       ;
  assign tx_phy_preflop_0 [  24] = 1'b0                       ;
  assign tx_phy_preflop_0 [  25] = 1'b0                       ;
  assign tx_phy_preflop_0 [  26] = 1'b0                       ;
  assign tx_phy_preflop_0 [  27] = 1'b0                       ;
  assign tx_phy_preflop_0 [  28] = 1'b0                       ;
  assign tx_phy_preflop_0 [  29] = 1'b0                       ;
  assign tx_phy_preflop_0 [  30] = 1'b0                       ;
  assign tx_phy_preflop_0 [  31] = 1'b0                       ;
  assign tx_phy_preflop_0 [  32] = 1'b0                       ;
  assign tx_phy_preflop_0 [  33] = 1'b0                       ;
  assign tx_phy_preflop_0 [  34] = 1'b0                       ;
  assign tx_phy_preflop_0 [  35] = 1'b0                       ;
  assign tx_phy_preflop_0 [  36] = 1'b0                       ;
  assign tx_phy_preflop_0 [  37] = 1'b0                       ;
  assign tx_phy_preflop_0 [  38] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [  39] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [  40] = 1'b0                       ;
  assign tx_phy_preflop_0 [  41] = 1'b0                       ;
  assign tx_phy_preflop_0 [  42] = 1'b0                       ;
  assign tx_phy_preflop_0 [  43] = 1'b0                       ;
  assign tx_phy_preflop_0 [  44] = 1'b0                       ;
  assign tx_phy_preflop_0 [  45] = 1'b0                       ;
  assign tx_phy_preflop_0 [  46] = 1'b0                       ;
  assign tx_phy_preflop_0 [  47] = 1'b0                       ;
  assign tx_phy_preflop_0 [  48] = 1'b0                       ;
  assign tx_phy_preflop_0 [  49] = 1'b0                       ;
  assign tx_phy_preflop_0 [  50] = 1'b0                       ;
  assign tx_phy_preflop_0 [  51] = 1'b0                       ;
  assign tx_phy_preflop_0 [  52] = 1'b0                       ;
  assign tx_phy_preflop_0 [  53] = 1'b0                       ;
  assign tx_phy_preflop_0 [  54] = 1'b0                       ;
  assign tx_phy_preflop_0 [  55] = 1'b0                       ;
  assign tx_phy_preflop_0 [  56] = 1'b0                       ;
  assign tx_phy_preflop_0 [  57] = 1'b0                       ;
  assign tx_phy_preflop_0 [  58] = 1'b0                       ;
  assign tx_phy_preflop_0 [  59] = 1'b0                       ;
  assign tx_phy_preflop_0 [  60] = 1'b0                       ;
  assign tx_phy_preflop_0 [  61] = 1'b0                       ;
  assign tx_phy_preflop_0 [  62] = 1'b0                       ;
  assign tx_phy_preflop_0 [  63] = 1'b0                       ;
  assign tx_phy_preflop_0 [  64] = 1'b0                       ;
  assign tx_phy_preflop_0 [  65] = 1'b0                       ;
  assign tx_phy_preflop_0 [  66] = 1'b0                       ;
  assign tx_phy_preflop_0 [  67] = 1'b0                       ;
  assign tx_phy_preflop_0 [  68] = 1'b0                       ;
  assign tx_phy_preflop_0 [  69] = 1'b0                       ;
  assign tx_phy_preflop_0 [  70] = 1'b0                       ;
  assign tx_phy_preflop_0 [  71] = 1'b0                       ;
  assign tx_phy_preflop_0 [  72] = 1'b0                       ;
  assign tx_phy_preflop_0 [  73] = 1'b0                       ;
  assign tx_phy_preflop_0 [  74] = 1'b0                       ;
  assign tx_phy_preflop_0 [  75] = 1'b0                       ;
  assign tx_phy_preflop_0 [  76] = 1'b0                       ;
  assign tx_phy_preflop_0 [  77] = 1'b0                       ;
  assign tx_phy_preflop_0 [  78] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [  79] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [   0] = tx_mrk_userbit[0]          ; // MARKER
  assign tx_phy_preflop_1 [   1] = tx_stb_userbit             ; // STROBE
  assign tx_phy_preflop_1 [   2] = 1'b0                       ;
  assign tx_phy_preflop_1 [   3] = 1'b0                       ;
  assign tx_phy_preflop_1 [   4] = 1'b0                       ;
  assign tx_phy_preflop_1 [   5] = 1'b0                       ;
  assign tx_phy_preflop_1 [   6] = 1'b0                       ;
  assign tx_phy_preflop_1 [   7] = 1'b0                       ;
  assign tx_phy_preflop_1 [   8] = 1'b0                       ;
  assign tx_phy_preflop_1 [   9] = 1'b0                       ;
  assign tx_phy_preflop_1 [  10] = 1'b0                       ;
  assign tx_phy_preflop_1 [  11] = 1'b0                       ;
  assign tx_phy_preflop_1 [  12] = 1'b0                       ;
  assign tx_phy_preflop_1 [  13] = 1'b0                       ;
  assign tx_phy_preflop_1 [  14] = 1'b0                       ;
  assign tx_phy_preflop_1 [  15] = 1'b0                       ;
  assign tx_phy_preflop_1 [  16] = 1'b0                       ;
  assign tx_phy_preflop_1 [  17] = 1'b0                       ;
  assign tx_phy_preflop_1 [  18] = 1'b0                       ;
  assign tx_phy_preflop_1 [  19] = 1'b0                       ;
  assign tx_phy_preflop_1 [  20] = 1'b0                       ;
  assign tx_phy_preflop_1 [  21] = 1'b0                       ;
  assign tx_phy_preflop_1 [  22] = 1'b0                       ;
  assign tx_phy_preflop_1 [  23] = 1'b0                       ;
  assign tx_phy_preflop_1 [  24] = 1'b0                       ;
  assign tx_phy_preflop_1 [  25] = 1'b0                       ;
  assign tx_phy_preflop_1 [  26] = 1'b0                       ;
  assign tx_phy_preflop_1 [  27] = 1'b0                       ;
  assign tx_phy_preflop_1 [  28] = 1'b0                       ;
  assign tx_phy_preflop_1 [  29] = 1'b0                       ;
  assign tx_phy_preflop_1 [  30] = 1'b0                       ;
  assign tx_phy_preflop_1 [  31] = 1'b0                       ;
  assign tx_phy_preflop_1 [  32] = 1'b0                       ;
  assign tx_phy_preflop_1 [  33] = 1'b0                       ;
  assign tx_phy_preflop_1 [  34] = 1'b0                       ;
  assign tx_phy_preflop_1 [  35] = 1'b0                       ;
  assign tx_phy_preflop_1 [  36] = 1'b0                       ;
  assign tx_phy_preflop_1 [  37] = 1'b0                       ;
  assign tx_phy_preflop_1 [  38] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [  39] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [  40] = 1'b0                       ;
  assign tx_phy_preflop_1 [  41] = 1'b0                       ;
  assign tx_phy_preflop_1 [  42] = 1'b0                       ;
  assign tx_phy_preflop_1 [  43] = 1'b0                       ;
  assign tx_phy_preflop_1 [  44] = 1'b0                       ;
  assign tx_phy_preflop_1 [  45] = 1'b0                       ;
  assign tx_phy_preflop_1 [  46] = 1'b0                       ;
  assign tx_phy_preflop_1 [  47] = 1'b0                       ;
  assign tx_phy_preflop_1 [  48] = 1'b0                       ;
  assign tx_phy_preflop_1 [  49] = 1'b0                       ;
  assign tx_phy_preflop_1 [  50] = 1'b0                       ;
  assign tx_phy_preflop_1 [  51] = 1'b0                       ;
  assign tx_phy_preflop_1 [  52] = 1'b0                       ;
  assign tx_phy_preflop_1 [  53] = 1'b0                       ;
  assign tx_phy_preflop_1 [  54] = 1'b0                       ;
  assign tx_phy_preflop_1 [  55] = 1'b0                       ;
  assign tx_phy_preflop_1 [  56] = 1'b0                       ;
  assign tx_phy_preflop_1 [  57] = 1'b0                       ;
  assign tx_phy_preflop_1 [  58] = 1'b0                       ;
  assign tx_phy_preflop_1 [  59] = 1'b0                       ;
  assign tx_phy_preflop_1 [  60] = 1'b0                       ;
  assign tx_phy_preflop_1 [  61] = 1'b0                       ;
  assign tx_phy_preflop_1 [  62] = 1'b0                       ;
  assign tx_phy_preflop_1 [  63] = 1'b0                       ;
  assign tx_phy_preflop_1 [  64] = 1'b0                       ;
  assign tx_phy_preflop_1 [  65] = 1'b0                       ;
  assign tx_phy_preflop_1 [  66] = 1'b0                       ;
  assign tx_phy_preflop_1 [  67] = 1'b0                       ;
  assign tx_phy_preflop_1 [  68] = 1'b0                       ;
  assign tx_phy_preflop_1 [  69] = 1'b0                       ;
  assign tx_phy_preflop_1 [  70] = 1'b0                       ;
  assign tx_phy_preflop_1 [  71] = 1'b0                       ;
  assign tx_phy_preflop_1 [  72] = 1'b0                       ;
  assign tx_phy_preflop_1 [  73] = 1'b0                       ;
  assign tx_phy_preflop_1 [  74] = 1'b0                       ;
  assign tx_phy_preflop_1 [  75] = 1'b0                       ;
  assign tx_phy_preflop_1 [  76] = 1'b0                       ;
  assign tx_phy_preflop_1 [  77] = 1'b0                       ;
  assign tx_phy_preflop_1 [  78] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [  79] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [  80] = tx_mrk_userbit[1]          ; // MARKER
  assign tx_phy_preflop_0 [  81] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_0 [  82] = tx_st_credit_r1            ;
  assign tx_phy_preflop_0 [  83] = 1'b0                       ;
  assign tx_phy_preflop_0 [  84] = 1'b0                       ;
  assign tx_phy_preflop_0 [  85] = 1'b0                       ;
  assign tx_phy_preflop_0 [  86] = 1'b0                       ;
  assign tx_phy_preflop_0 [  87] = 1'b0                       ;
  assign tx_phy_preflop_0 [  88] = 1'b0                       ;
  assign tx_phy_preflop_0 [  89] = 1'b0                       ;
  assign tx_phy_preflop_0 [  90] = 1'b0                       ;
  assign tx_phy_preflop_0 [  91] = 1'b0                       ;
  assign tx_phy_preflop_0 [  92] = 1'b0                       ;
  assign tx_phy_preflop_0 [  93] = 1'b0                       ;
  assign tx_phy_preflop_0 [  94] = 1'b0                       ;
  assign tx_phy_preflop_0 [  95] = 1'b0                       ;
  assign tx_phy_preflop_0 [  96] = 1'b0                       ;
  assign tx_phy_preflop_0 [  97] = 1'b0                       ;
  assign tx_phy_preflop_0 [  98] = 1'b0                       ;
  assign tx_phy_preflop_0 [  99] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 100] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 101] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 102] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 103] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 104] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 105] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 106] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 107] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 108] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 109] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 110] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 111] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 112] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 113] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 114] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 115] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 116] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 117] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 118] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 119] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 120] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 121] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 122] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 123] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 124] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 125] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 126] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 127] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 128] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 129] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 130] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 131] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 132] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 133] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 134] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 135] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 136] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 137] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 138] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 139] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 140] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 141] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 142] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 143] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 144] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 145] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 146] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 147] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 148] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 149] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 150] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 151] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 152] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 153] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 154] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 155] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 156] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 157] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 158] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 159] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [  80] = tx_mrk_userbit[1]          ; // MARKER
  assign tx_phy_preflop_1 [  81] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_1 [  82] = 1'b0                       ;
  assign tx_phy_preflop_1 [  83] = 1'b0                       ;
  assign tx_phy_preflop_1 [  84] = 1'b0                       ;
  assign tx_phy_preflop_1 [  85] = 1'b0                       ;
  assign tx_phy_preflop_1 [  86] = 1'b0                       ;
  assign tx_phy_preflop_1 [  87] = 1'b0                       ;
  assign tx_phy_preflop_1 [  88] = 1'b0                       ;
  assign tx_phy_preflop_1 [  89] = 1'b0                       ;
  assign tx_phy_preflop_1 [  90] = 1'b0                       ;
  assign tx_phy_preflop_1 [  91] = 1'b0                       ;
  assign tx_phy_preflop_1 [  92] = 1'b0                       ;
  assign tx_phy_preflop_1 [  93] = 1'b0                       ;
  assign tx_phy_preflop_1 [  94] = 1'b0                       ;
  assign tx_phy_preflop_1 [  95] = 1'b0                       ;
  assign tx_phy_preflop_1 [  96] = 1'b0                       ;
  assign tx_phy_preflop_1 [  97] = 1'b0                       ;
  assign tx_phy_preflop_1 [  98] = 1'b0                       ;
  assign tx_phy_preflop_1 [  99] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 100] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 101] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 102] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 103] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 104] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 105] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 106] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 107] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 108] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 109] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 110] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 111] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 112] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 113] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 114] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 115] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 116] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 117] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 118] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 119] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 120] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 121] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 122] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 123] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 124] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 125] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 126] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 127] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 128] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 129] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 130] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 131] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 132] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 133] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 134] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 135] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 136] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 137] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 138] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 139] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 140] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 141] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 142] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 143] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 144] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 145] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 146] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 147] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 148] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 149] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 150] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 151] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 152] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 153] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 154] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 155] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 156] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 157] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 158] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 159] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 160] = tx_mrk_userbit[2]          ; // MARKER
  assign tx_phy_preflop_0 [ 161] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_0 [ 162] = tx_st_credit_r2            ;
  assign tx_phy_preflop_0 [ 163] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 164] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 165] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 166] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 167] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 168] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 169] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 170] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 171] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 172] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 173] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 174] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 175] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 176] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 177] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 178] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 179] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 180] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 181] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 182] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 183] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 184] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 185] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 186] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 187] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 188] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 189] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 190] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 191] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 192] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 193] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 194] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 195] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 196] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 197] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 198] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 199] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 200] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 201] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 202] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 203] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 204] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 205] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 206] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 207] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 208] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 209] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 210] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 211] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 212] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 213] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 214] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 215] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 216] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 217] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 218] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 219] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 220] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 221] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 222] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 223] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 224] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 225] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 226] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 227] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 228] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 229] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 230] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 231] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 232] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 233] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 234] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 235] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 236] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 237] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 238] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 239] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 160] = tx_mrk_userbit[2]          ; // MARKER
  assign tx_phy_preflop_1 [ 161] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_1 [ 162] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 163] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 164] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 165] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 166] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 167] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 168] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 169] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 170] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 171] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 172] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 173] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 174] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 175] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 176] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 177] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 178] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 179] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 180] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 181] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 182] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 183] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 184] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 185] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 186] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 187] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 188] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 189] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 190] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 191] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 192] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 193] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 194] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 195] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 196] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 197] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 198] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 199] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 200] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 201] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 202] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 203] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 204] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 205] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 206] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 207] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 208] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 209] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 210] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 211] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 212] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 213] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 214] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 215] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 216] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 217] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 218] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 219] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 220] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 221] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 222] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 223] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 224] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 225] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 226] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 227] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 228] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 229] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 230] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 231] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 232] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 233] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 234] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 235] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 236] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 237] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 238] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 239] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 240] = tx_mrk_userbit[3]          ; // MARKER
  assign tx_phy_preflop_0 [ 241] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_0 [ 242] = tx_st_credit_r3            ;
  assign tx_phy_preflop_0 [ 243] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 244] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 245] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 246] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 247] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 248] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 249] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 250] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 251] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 252] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 253] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 254] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 255] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 256] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 257] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 258] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 259] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 260] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 261] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 262] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 263] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 264] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 265] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 266] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 267] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 268] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 269] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 270] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 271] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 272] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 273] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 274] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 275] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 276] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 277] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 278] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 279] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 280] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 281] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 282] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 283] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 284] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 285] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 286] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 287] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 288] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 289] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 290] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 291] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 292] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 293] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 294] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 295] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 296] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 297] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 298] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 299] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 300] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 301] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 302] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 303] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 304] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 305] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 306] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 307] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 308] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 309] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 310] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 311] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 312] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 313] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 314] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 315] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 316] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 317] = 1'b0                       ;
  assign tx_phy_preflop_0 [ 318] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 319] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 240] = tx_mrk_userbit[3]          ; // MARKER
  assign tx_phy_preflop_1 [ 241] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_1 [ 242] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 243] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 244] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 245] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 246] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 247] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 248] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 249] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 250] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 251] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 252] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 253] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 254] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 255] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 256] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 257] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 258] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 259] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 260] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 261] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 262] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 263] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 264] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 265] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 266] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 267] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 268] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 269] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 270] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 271] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 272] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 273] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 274] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 275] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 276] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 277] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 278] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 279] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 280] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 281] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 282] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 283] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 284] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 285] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 286] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 287] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 288] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 289] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 290] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 291] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 292] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 293] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 294] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 295] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 296] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 297] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 298] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 299] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 300] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 301] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 302] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 303] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 304] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 305] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 306] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 307] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 308] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 309] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 310] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 311] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 312] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 313] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 314] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 315] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 316] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 317] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 318] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 319] = 1'b0                       ; // DBI
// TX Section
//////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////
// RX Section

//   RX_CH_WIDTH           = 320; // Gen2Only running at Quarter Rate
//   RX_DATA_WIDTH         = 296; // Usable Data per Channel
//   RX_PERSISTENT_STROBE  = 1'b1;
//   RX_PERSISTENT_MARKER  = 1'b1;
//   RX_STROBE_GEN2_LOC    = 'd1;
//   RX_MARKER_GEN2_LOC    = 'd0;
//   RX_STROBE_GEN1_LOC    = 'd38;
//   RX_MARKER_GEN1_LOC    = 'd39;
//   RX_ENABLE_STROBE      = 1'b1;
//   RX_ENABLE_MARKER      = 1'b1;
//   RX_DBI_PRESENT        = 1'b1;
//   RX_REG_PHY            = 1'b0;

  localparam RX_REG_PHY    = 1'b0;  // If set, this enables boundary FF for timing reasons

  logic [ 319:   0]                              rx_phy_postflop_0             ;
  logic [ 319:   0]                              rx_phy_postflop_1             ;
  logic [ 319:   0]                              rx_phy_flop_0_reg             ;
  logic [ 319:   0]                              rx_phy_flop_1_reg             ;

  always_ff @(posedge clk_rd or negedge rst_rd_n)
  if (~rst_rd_n)
  begin
    rx_phy_flop_0_reg                       <= 320'b0                                  ;
    rx_phy_flop_1_reg                       <= 320'b0                                  ;
  end
  else
  begin
    rx_phy_flop_0_reg                       <= rx_phy0                                 ;
    rx_phy_flop_1_reg                       <= rx_phy1                                 ;
  end


  assign rx_phy_postflop_0                  = RX_REG_PHY ? rx_phy_flop_0_reg : rx_phy0               ;
  assign rx_phy_postflop_1                  = RX_REG_PHY ? rx_phy_flop_1_reg : rx_phy1               ;

  logic                                          rx_st_pushbit_r0              ;
  logic                                          rx_st_pushbit_r1              ;
  logic                                          rx_st_pushbit_r2              ;
  logic                                          rx_st_pushbit_r3              ;

  assign rx_st_pushbit        = rx_st_pushbit_r0    |
                                rx_st_pushbit_r1    |
                                rx_st_pushbit_r2    |
                                rx_st_pushbit_r3    ;

//       MARKER                     = rx_phy_postflop_0 [   0]
//       STROBE                     = rx_phy_postflop_0 [   1]
  assign rx_st_pushbit_r0           = rx_phy_postflop_0 [   2];
  assign rx_st_data          [   0] = rx_phy_postflop_0 [   3];
  assign rx_st_data          [   1] = rx_phy_postflop_0 [   4];
  assign rx_st_data          [   2] = rx_phy_postflop_0 [   5];
  assign rx_st_data          [   3] = rx_phy_postflop_0 [   6];
  assign rx_st_data          [   4] = rx_phy_postflop_0 [   7];
  assign rx_st_data          [   5] = rx_phy_postflop_0 [   8];
  assign rx_st_data          [   6] = rx_phy_postflop_0 [   9];
  assign rx_st_data          [   7] = rx_phy_postflop_0 [  10];
  assign rx_st_data          [   8] = rx_phy_postflop_0 [  11];
  assign rx_st_data          [   9] = rx_phy_postflop_0 [  12];
  assign rx_st_data          [  10] = rx_phy_postflop_0 [  13];
  assign rx_st_data          [  11] = rx_phy_postflop_0 [  14];
  assign rx_st_data          [  12] = rx_phy_postflop_0 [  15];
  assign rx_st_data          [  13] = rx_phy_postflop_0 [  16];
  assign rx_st_data          [  14] = rx_phy_postflop_0 [  17];
  assign rx_st_data          [  15] = rx_phy_postflop_0 [  18];
  assign rx_st_data          [  16] = rx_phy_postflop_0 [  19];
  assign rx_st_data          [  17] = rx_phy_postflop_0 [  20];
  assign rx_st_data          [  18] = rx_phy_postflop_0 [  21];
  assign rx_st_data          [  19] = rx_phy_postflop_0 [  22];
  assign rx_st_data          [  20] = rx_phy_postflop_0 [  23];
  assign rx_st_data          [  21] = rx_phy_postflop_0 [  24];
  assign rx_st_data          [  22] = rx_phy_postflop_0 [  25];
  assign rx_st_data          [  23] = rx_phy_postflop_0 [  26];
  assign rx_st_data          [  24] = rx_phy_postflop_0 [  27];
  assign rx_st_data          [  25] = rx_phy_postflop_0 [  28];
  assign rx_st_data          [  26] = rx_phy_postflop_0 [  29];
  assign rx_st_data          [  27] = rx_phy_postflop_0 [  30];
  assign rx_st_data          [  28] = rx_phy_postflop_0 [  31];
  assign rx_st_data          [  29] = rx_phy_postflop_0 [  32];
  assign rx_st_data          [  30] = rx_phy_postflop_0 [  33];
  assign rx_st_data          [  31] = rx_phy_postflop_0 [  34];
  assign rx_st_data          [  32] = rx_phy_postflop_0 [  35];
  assign rx_st_data          [  33] = rx_phy_postflop_0 [  36];
  assign rx_st_data          [  34] = rx_phy_postflop_0 [  37];
//       DBI                        = rx_phy_postflop_0 [  38];
//       DBI                        = rx_phy_postflop_0 [  39];
  assign rx_st_data          [  35] = rx_phy_postflop_0 [  40];
  assign rx_st_data          [  36] = rx_phy_postflop_0 [  41];
  assign rx_st_data          [  37] = rx_phy_postflop_0 [  42];
  assign rx_st_data          [  38] = rx_phy_postflop_0 [  43];
  assign rx_st_data          [  39] = rx_phy_postflop_0 [  44];
  assign rx_st_data          [  40] = rx_phy_postflop_0 [  45];
  assign rx_st_data          [  41] = rx_phy_postflop_0 [  46];
  assign rx_st_data          [  42] = rx_phy_postflop_0 [  47];
  assign rx_st_data          [  43] = rx_phy_postflop_0 [  48];
  assign rx_st_data          [  44] = rx_phy_postflop_0 [  49];
  assign rx_st_data          [  45] = rx_phy_postflop_0 [  50];
  assign rx_st_data          [  46] = rx_phy_postflop_0 [  51];
  assign rx_st_data          [  47] = rx_phy_postflop_0 [  52];
  assign rx_st_data          [  48] = rx_phy_postflop_0 [  53];
  assign rx_st_data          [  49] = rx_phy_postflop_0 [  54];
  assign rx_st_data          [  50] = rx_phy_postflop_0 [  55];
  assign rx_st_data          [  51] = rx_phy_postflop_0 [  56];
  assign rx_st_data          [  52] = rx_phy_postflop_0 [  57];
  assign rx_st_data          [  53] = rx_phy_postflop_0 [  58];
  assign rx_st_data          [  54] = rx_phy_postflop_0 [  59];
  assign rx_st_data          [  55] = rx_phy_postflop_0 [  60];
  assign rx_st_data          [  56] = rx_phy_postflop_0 [  61];
  assign rx_st_data          [  57] = rx_phy_postflop_0 [  62];
  assign rx_st_data          [  58] = rx_phy_postflop_0 [  63];
  assign rx_st_data          [  59] = rx_phy_postflop_0 [  64];
  assign rx_st_data          [  60] = rx_phy_postflop_0 [  65];
  assign rx_st_data          [  61] = rx_phy_postflop_0 [  66];
  assign rx_st_data          [  62] = rx_phy_postflop_0 [  67];
  assign rx_st_data          [  63] = rx_phy_postflop_0 [  68];
  assign rx_st_data          [  64] = rx_phy_postflop_0 [  69];
  assign rx_st_data          [  65] = rx_phy_postflop_0 [  70];
  assign rx_st_data          [  66] = rx_phy_postflop_0 [  71];
  assign rx_st_data          [  67] = rx_phy_postflop_0 [  72];
  assign rx_st_data          [  68] = rx_phy_postflop_0 [  73];
  assign rx_st_data          [  69] = rx_phy_postflop_0 [  74];
  assign rx_st_data          [  70] = rx_phy_postflop_0 [  75];
  assign rx_st_data          [  71] = rx_phy_postflop_0 [  76];
  assign rx_st_data          [  72] = rx_phy_postflop_0 [  77];
//       DBI                        = rx_phy_postflop_0 [  78];
//       DBI                        = rx_phy_postflop_0 [  79];
//       MARKER                     = rx_phy_postflop_1 [   0]
//       STROBE                     = rx_phy_postflop_1 [   1]
  assign rx_st_data          [  73] = rx_phy_postflop_1 [   2];
  assign rx_st_data          [  74] = rx_phy_postflop_1 [   3];
  assign rx_st_data          [  75] = rx_phy_postflop_1 [   4];
  assign rx_st_data          [  76] = rx_phy_postflop_1 [   5];
  assign rx_st_data          [  77] = rx_phy_postflop_1 [   6];
  assign rx_st_data          [  78] = rx_phy_postflop_1 [   7];
  assign rx_st_data          [  79] = rx_phy_postflop_1 [   8];
  assign rx_st_data          [  80] = rx_phy_postflop_1 [   9];
  assign rx_st_data          [  81] = rx_phy_postflop_1 [  10];
  assign rx_st_data          [  82] = rx_phy_postflop_1 [  11];
  assign rx_st_data          [  83] = rx_phy_postflop_1 [  12];
  assign rx_st_data          [  84] = rx_phy_postflop_1 [  13];
  assign rx_st_data          [  85] = rx_phy_postflop_1 [  14];
  assign rx_st_data          [  86] = rx_phy_postflop_1 [  15];
  assign rx_st_data          [  87] = rx_phy_postflop_1 [  16];
  assign rx_st_data          [  88] = rx_phy_postflop_1 [  17];
  assign rx_st_data          [  89] = rx_phy_postflop_1 [  18];
  assign rx_st_data          [  90] = rx_phy_postflop_1 [  19];
  assign rx_st_data          [  91] = rx_phy_postflop_1 [  20];
  assign rx_st_data          [  92] = rx_phy_postflop_1 [  21];
  assign rx_st_data          [  93] = rx_phy_postflop_1 [  22];
  assign rx_st_data          [  94] = rx_phy_postflop_1 [  23];
  assign rx_st_data          [  95] = rx_phy_postflop_1 [  24];
  assign rx_st_data          [  96] = rx_phy_postflop_1 [  25];
  assign rx_st_data          [  97] = rx_phy_postflop_1 [  26];
  assign rx_st_data          [  98] = rx_phy_postflop_1 [  27];
  assign rx_st_data          [  99] = rx_phy_postflop_1 [  28];
  assign rx_st_data          [ 100] = rx_phy_postflop_1 [  29];
  assign rx_st_data          [ 101] = rx_phy_postflop_1 [  30];
  assign rx_st_data          [ 102] = rx_phy_postflop_1 [  31];
  assign rx_st_data          [ 103] = rx_phy_postflop_1 [  32];
  assign rx_st_data          [ 104] = rx_phy_postflop_1 [  33];
  assign rx_st_data          [ 105] = rx_phy_postflop_1 [  34];
  assign rx_st_data          [ 106] = rx_phy_postflop_1 [  35];
  assign rx_st_data          [ 107] = rx_phy_postflop_1 [  36];
  assign rx_st_data          [ 108] = rx_phy_postflop_1 [  37];
//       DBI                        = rx_phy_postflop_1 [  38];
//       DBI                        = rx_phy_postflop_1 [  39];
  assign rx_st_data          [ 109] = rx_phy_postflop_1 [  40];
  assign rx_st_data          [ 110] = rx_phy_postflop_1 [  41];
  assign rx_st_data          [ 111] = rx_phy_postflop_1 [  42];
  assign rx_st_data          [ 112] = rx_phy_postflop_1 [  43];
  assign rx_st_data          [ 113] = rx_phy_postflop_1 [  44];
  assign rx_st_data          [ 114] = rx_phy_postflop_1 [  45];
  assign rx_st_data          [ 115] = rx_phy_postflop_1 [  46];
  assign rx_st_data          [ 116] = rx_phy_postflop_1 [  47];
  assign rx_st_data          [ 117] = rx_phy_postflop_1 [  48];
  assign rx_st_data          [ 118] = rx_phy_postflop_1 [  49];
  assign rx_st_data          [ 119] = rx_phy_postflop_1 [  50];
  assign rx_st_data          [ 120] = rx_phy_postflop_1 [  51];
  assign rx_st_data          [ 121] = rx_phy_postflop_1 [  52];
  assign rx_st_data          [ 122] = rx_phy_postflop_1 [  53];
  assign rx_st_data          [ 123] = rx_phy_postflop_1 [  54];
  assign rx_st_data          [ 124] = rx_phy_postflop_1 [  55];
  assign rx_st_data          [ 125] = rx_phy_postflop_1 [  56];
  assign rx_st_data          [ 126] = rx_phy_postflop_1 [  57];
  assign rx_st_data          [ 127] = rx_phy_postflop_1 [  58];
  assign rx_st_data          [ 128] = rx_phy_postflop_1 [  59];
  assign rx_st_data          [ 129] = rx_phy_postflop_1 [  60];
  assign rx_st_data          [ 130] = rx_phy_postflop_1 [  61];
  assign rx_st_data          [ 131] = rx_phy_postflop_1 [  62];
  assign rx_st_data          [ 132] = rx_phy_postflop_1 [  63];
  assign rx_st_data          [ 133] = rx_phy_postflop_1 [  64];
  assign rx_st_data          [ 134] = rx_phy_postflop_1 [  65];
  assign rx_st_data          [ 135] = rx_phy_postflop_1 [  66];
  assign rx_st_data          [ 136] = rx_phy_postflop_1 [  67];
  assign rx_st_data          [ 137] = rx_phy_postflop_1 [  68];
  assign rx_st_data          [ 138] = rx_phy_postflop_1 [  69];
  assign rx_st_data          [ 139] = rx_phy_postflop_1 [  70];
  assign rx_st_data          [ 140] = rx_phy_postflop_1 [  71];
  assign rx_st_data          [ 141] = rx_phy_postflop_1 [  72];
  assign rx_st_data          [ 142] = rx_phy_postflop_1 [  73];
  assign rx_st_data          [ 143] = rx_phy_postflop_1 [  74];
  assign rx_st_data          [ 144] = rx_phy_postflop_1 [  75];
//       nc                         = rx_phy_postflop_1 [  76];
//       nc                         = rx_phy_postflop_1 [  77];
//       DBI                        = rx_phy_postflop_1 [  78];
//       DBI                        = rx_phy_postflop_1 [  79];
//       MARKER                     = rx_phy_postflop_0 [  80]
//       STROBE                     = rx_phy_postflop_0 [  81]
  assign rx_st_pushbit_r1           = rx_phy_postflop_0 [  82];
  assign rx_st_data          [ 145] = rx_phy_postflop_0 [  83];
  assign rx_st_data          [ 146] = rx_phy_postflop_0 [  84];
  assign rx_st_data          [ 147] = rx_phy_postflop_0 [  85];
  assign rx_st_data          [ 148] = rx_phy_postflop_0 [  86];
  assign rx_st_data          [ 149] = rx_phy_postflop_0 [  87];
  assign rx_st_data          [ 150] = rx_phy_postflop_0 [  88];
  assign rx_st_data          [ 151] = rx_phy_postflop_0 [  89];
  assign rx_st_data          [ 152] = rx_phy_postflop_0 [  90];
  assign rx_st_data          [ 153] = rx_phy_postflop_0 [  91];
  assign rx_st_data          [ 154] = rx_phy_postflop_0 [  92];
  assign rx_st_data          [ 155] = rx_phy_postflop_0 [  93];
  assign rx_st_data          [ 156] = rx_phy_postflop_0 [  94];
  assign rx_st_data          [ 157] = rx_phy_postflop_0 [  95];
  assign rx_st_data          [ 158] = rx_phy_postflop_0 [  96];
  assign rx_st_data          [ 159] = rx_phy_postflop_0 [  97];
  assign rx_st_data          [ 160] = rx_phy_postflop_0 [  98];
  assign rx_st_data          [ 161] = rx_phy_postflop_0 [  99];
  assign rx_st_data          [ 162] = rx_phy_postflop_0 [ 100];
  assign rx_st_data          [ 163] = rx_phy_postflop_0 [ 101];
  assign rx_st_data          [ 164] = rx_phy_postflop_0 [ 102];
  assign rx_st_data          [ 165] = rx_phy_postflop_0 [ 103];
  assign rx_st_data          [ 166] = rx_phy_postflop_0 [ 104];
  assign rx_st_data          [ 167] = rx_phy_postflop_0 [ 105];
  assign rx_st_data          [ 168] = rx_phy_postflop_0 [ 106];
  assign rx_st_data          [ 169] = rx_phy_postflop_0 [ 107];
  assign rx_st_data          [ 170] = rx_phy_postflop_0 [ 108];
  assign rx_st_data          [ 171] = rx_phy_postflop_0 [ 109];
  assign rx_st_data          [ 172] = rx_phy_postflop_0 [ 110];
  assign rx_st_data          [ 173] = rx_phy_postflop_0 [ 111];
  assign rx_st_data          [ 174] = rx_phy_postflop_0 [ 112];
  assign rx_st_data          [ 175] = rx_phy_postflop_0 [ 113];
  assign rx_st_data          [ 176] = rx_phy_postflop_0 [ 114];
  assign rx_st_data          [ 177] = rx_phy_postflop_0 [ 115];
  assign rx_st_data          [ 178] = rx_phy_postflop_0 [ 116];
  assign rx_st_data          [ 179] = rx_phy_postflop_0 [ 117];
//       DBI                        = rx_phy_postflop_0 [ 118];
//       DBI                        = rx_phy_postflop_0 [ 119];
  assign rx_st_data          [ 180] = rx_phy_postflop_0 [ 120];
  assign rx_st_data          [ 181] = rx_phy_postflop_0 [ 121];
  assign rx_st_data          [ 182] = rx_phy_postflop_0 [ 122];
  assign rx_st_data          [ 183] = rx_phy_postflop_0 [ 123];
  assign rx_st_data          [ 184] = rx_phy_postflop_0 [ 124];
  assign rx_st_data          [ 185] = rx_phy_postflop_0 [ 125];
  assign rx_st_data          [ 186] = rx_phy_postflop_0 [ 126];
  assign rx_st_data          [ 187] = rx_phy_postflop_0 [ 127];
  assign rx_st_data          [ 188] = rx_phy_postflop_0 [ 128];
  assign rx_st_data          [ 189] = rx_phy_postflop_0 [ 129];
  assign rx_st_data          [ 190] = rx_phy_postflop_0 [ 130];
  assign rx_st_data          [ 191] = rx_phy_postflop_0 [ 131];
  assign rx_st_data          [ 192] = rx_phy_postflop_0 [ 132];
  assign rx_st_data          [ 193] = rx_phy_postflop_0 [ 133];
  assign rx_st_data          [ 194] = rx_phy_postflop_0 [ 134];
  assign rx_st_data          [ 195] = rx_phy_postflop_0 [ 135];
  assign rx_st_data          [ 196] = rx_phy_postflop_0 [ 136];
  assign rx_st_data          [ 197] = rx_phy_postflop_0 [ 137];
  assign rx_st_data          [ 198] = rx_phy_postflop_0 [ 138];
  assign rx_st_data          [ 199] = rx_phy_postflop_0 [ 139];
  assign rx_st_data          [ 200] = rx_phy_postflop_0 [ 140];
  assign rx_st_data          [ 201] = rx_phy_postflop_0 [ 141];
  assign rx_st_data          [ 202] = rx_phy_postflop_0 [ 142];
  assign rx_st_data          [ 203] = rx_phy_postflop_0 [ 143];
  assign rx_st_data          [ 204] = rx_phy_postflop_0 [ 144];
  assign rx_st_data          [ 205] = rx_phy_postflop_0 [ 145];
  assign rx_st_data          [ 206] = rx_phy_postflop_0 [ 146];
  assign rx_st_data          [ 207] = rx_phy_postflop_0 [ 147];
  assign rx_st_data          [ 208] = rx_phy_postflop_0 [ 148];
  assign rx_st_data          [ 209] = rx_phy_postflop_0 [ 149];
  assign rx_st_data          [ 210] = rx_phy_postflop_0 [ 150];
  assign rx_st_data          [ 211] = rx_phy_postflop_0 [ 151];
  assign rx_st_data          [ 212] = rx_phy_postflop_0 [ 152];
  assign rx_st_data          [ 213] = rx_phy_postflop_0 [ 153];
  assign rx_st_data          [ 214] = rx_phy_postflop_0 [ 154];
  assign rx_st_data          [ 215] = rx_phy_postflop_0 [ 155];
  assign rx_st_data          [ 216] = rx_phy_postflop_0 [ 156];
  assign rx_st_data          [ 217] = rx_phy_postflop_0 [ 157];
//       DBI                        = rx_phy_postflop_0 [ 158];
//       DBI                        = rx_phy_postflop_0 [ 159];
//       MARKER                     = rx_phy_postflop_1 [  80]
//       STROBE                     = rx_phy_postflop_1 [  81]
  assign rx_st_data          [ 218] = rx_phy_postflop_1 [  82];
  assign rx_st_data          [ 219] = rx_phy_postflop_1 [  83];
  assign rx_st_data          [ 220] = rx_phy_postflop_1 [  84];
  assign rx_st_data          [ 221] = rx_phy_postflop_1 [  85];
  assign rx_st_data          [ 222] = rx_phy_postflop_1 [  86];
  assign rx_st_data          [ 223] = rx_phy_postflop_1 [  87];
  assign rx_st_data          [ 224] = rx_phy_postflop_1 [  88];
  assign rx_st_data          [ 225] = rx_phy_postflop_1 [  89];
  assign rx_st_data          [ 226] = rx_phy_postflop_1 [  90];
  assign rx_st_data          [ 227] = rx_phy_postflop_1 [  91];
  assign rx_st_data          [ 228] = rx_phy_postflop_1 [  92];
  assign rx_st_data          [ 229] = rx_phy_postflop_1 [  93];
  assign rx_st_data          [ 230] = rx_phy_postflop_1 [  94];
  assign rx_st_data          [ 231] = rx_phy_postflop_1 [  95];
  assign rx_st_data          [ 232] = rx_phy_postflop_1 [  96];
  assign rx_st_data          [ 233] = rx_phy_postflop_1 [  97];
  assign rx_st_data          [ 234] = rx_phy_postflop_1 [  98];
  assign rx_st_data          [ 235] = rx_phy_postflop_1 [  99];
  assign rx_st_data          [ 236] = rx_phy_postflop_1 [ 100];
  assign rx_st_data          [ 237] = rx_phy_postflop_1 [ 101];
  assign rx_st_data          [ 238] = rx_phy_postflop_1 [ 102];
  assign rx_st_data          [ 239] = rx_phy_postflop_1 [ 103];
  assign rx_st_data          [ 240] = rx_phy_postflop_1 [ 104];
  assign rx_st_data          [ 241] = rx_phy_postflop_1 [ 105];
  assign rx_st_data          [ 242] = rx_phy_postflop_1 [ 106];
  assign rx_st_data          [ 243] = rx_phy_postflop_1 [ 107];
  assign rx_st_data          [ 244] = rx_phy_postflop_1 [ 108];
  assign rx_st_data          [ 245] = rx_phy_postflop_1 [ 109];
  assign rx_st_data          [ 246] = rx_phy_postflop_1 [ 110];
  assign rx_st_data          [ 247] = rx_phy_postflop_1 [ 111];
  assign rx_st_data          [ 248] = rx_phy_postflop_1 [ 112];
  assign rx_st_data          [ 249] = rx_phy_postflop_1 [ 113];
  assign rx_st_data          [ 250] = rx_phy_postflop_1 [ 114];
  assign rx_st_data          [ 251] = rx_phy_postflop_1 [ 115];
  assign rx_st_data          [ 252] = rx_phy_postflop_1 [ 116];
  assign rx_st_data          [ 253] = rx_phy_postflop_1 [ 117];
//       DBI                        = rx_phy_postflop_1 [ 118];
//       DBI                        = rx_phy_postflop_1 [ 119];
  assign rx_st_data          [ 254] = rx_phy_postflop_1 [ 120];
  assign rx_st_data          [ 255] = rx_phy_postflop_1 [ 121];
  assign rx_st_data          [ 256] = rx_phy_postflop_1 [ 122];
  assign rx_st_data          [ 257] = rx_phy_postflop_1 [ 123];
  assign rx_st_data          [ 258] = rx_phy_postflop_1 [ 124];
  assign rx_st_data          [ 259] = rx_phy_postflop_1 [ 125];
  assign rx_st_data          [ 260] = rx_phy_postflop_1 [ 126];
  assign rx_st_data          [ 261] = rx_phy_postflop_1 [ 127];
  assign rx_st_data          [ 262] = rx_phy_postflop_1 [ 128];
  assign rx_st_data          [ 263] = rx_phy_postflop_1 [ 129];
  assign rx_st_data          [ 264] = rx_phy_postflop_1 [ 130];
  assign rx_st_data          [ 265] = rx_phy_postflop_1 [ 131];
  assign rx_st_data          [ 266] = rx_phy_postflop_1 [ 132];
  assign rx_st_data          [ 267] = rx_phy_postflop_1 [ 133];
  assign rx_st_data          [ 268] = rx_phy_postflop_1 [ 134];
  assign rx_st_data          [ 269] = rx_phy_postflop_1 [ 135];
  assign rx_st_data          [ 270] = rx_phy_postflop_1 [ 136];
  assign rx_st_data          [ 271] = rx_phy_postflop_1 [ 137];
  assign rx_st_data          [ 272] = rx_phy_postflop_1 [ 138];
  assign rx_st_data          [ 273] = rx_phy_postflop_1 [ 139];
  assign rx_st_data          [ 274] = rx_phy_postflop_1 [ 140];
  assign rx_st_data          [ 275] = rx_phy_postflop_1 [ 141];
  assign rx_st_data          [ 276] = rx_phy_postflop_1 [ 142];
  assign rx_st_data          [ 277] = rx_phy_postflop_1 [ 143];
  assign rx_st_data          [ 278] = rx_phy_postflop_1 [ 144];
  assign rx_st_data          [ 279] = rx_phy_postflop_1 [ 145];
  assign rx_st_data          [ 280] = rx_phy_postflop_1 [ 146];
  assign rx_st_data          [ 281] = rx_phy_postflop_1 [ 147];
  assign rx_st_data          [ 282] = rx_phy_postflop_1 [ 148];
  assign rx_st_data          [ 283] = rx_phy_postflop_1 [ 149];
  assign rx_st_data          [ 284] = rx_phy_postflop_1 [ 150];
  assign rx_st_data          [ 285] = rx_phy_postflop_1 [ 151];
  assign rx_st_data          [ 286] = rx_phy_postflop_1 [ 152];
  assign rx_st_data          [ 287] = rx_phy_postflop_1 [ 153];
  assign rx_st_data          [ 288] = rx_phy_postflop_1 [ 154];
  assign rx_st_data          [ 289] = rx_phy_postflop_1 [ 155];
//       nc                         = rx_phy_postflop_1 [ 156];
//       nc                         = rx_phy_postflop_1 [ 157];
//       DBI                        = rx_phy_postflop_1 [ 158];
//       DBI                        = rx_phy_postflop_1 [ 159];
//       MARKER                     = rx_phy_postflop_0 [ 160]
//       STROBE                     = rx_phy_postflop_0 [ 161]
  assign rx_st_pushbit_r2           = rx_phy_postflop_0 [ 162];
  assign rx_st_data          [ 290] = rx_phy_postflop_0 [ 163];
  assign rx_st_data          [ 291] = rx_phy_postflop_0 [ 164];
  assign rx_st_data          [ 292] = rx_phy_postflop_0 [ 165];
  assign rx_st_data          [ 293] = rx_phy_postflop_0 [ 166];
  assign rx_st_data          [ 294] = rx_phy_postflop_0 [ 167];
  assign rx_st_data          [ 295] = rx_phy_postflop_0 [ 168];
  assign rx_st_data          [ 296] = rx_phy_postflop_0 [ 169];
  assign rx_st_data          [ 297] = rx_phy_postflop_0 [ 170];
  assign rx_st_data          [ 298] = rx_phy_postflop_0 [ 171];
  assign rx_st_data          [ 299] = rx_phy_postflop_0 [ 172];
  assign rx_st_data          [ 300] = rx_phy_postflop_0 [ 173];
  assign rx_st_data          [ 301] = rx_phy_postflop_0 [ 174];
  assign rx_st_data          [ 302] = rx_phy_postflop_0 [ 175];
  assign rx_st_data          [ 303] = rx_phy_postflop_0 [ 176];
  assign rx_st_data          [ 304] = rx_phy_postflop_0 [ 177];
  assign rx_st_data          [ 305] = rx_phy_postflop_0 [ 178];
  assign rx_st_data          [ 306] = rx_phy_postflop_0 [ 179];
  assign rx_st_data          [ 307] = rx_phy_postflop_0 [ 180];
  assign rx_st_data          [ 308] = rx_phy_postflop_0 [ 181];
  assign rx_st_data          [ 309] = rx_phy_postflop_0 [ 182];
  assign rx_st_data          [ 310] = rx_phy_postflop_0 [ 183];
  assign rx_st_data          [ 311] = rx_phy_postflop_0 [ 184];
  assign rx_st_data          [ 312] = rx_phy_postflop_0 [ 185];
  assign rx_st_data          [ 313] = rx_phy_postflop_0 [ 186];
  assign rx_st_data          [ 314] = rx_phy_postflop_0 [ 187];
  assign rx_st_data          [ 315] = rx_phy_postflop_0 [ 188];
  assign rx_st_data          [ 316] = rx_phy_postflop_0 [ 189];
  assign rx_st_data          [ 317] = rx_phy_postflop_0 [ 190];
  assign rx_st_data          [ 318] = rx_phy_postflop_0 [ 191];
  assign rx_st_data          [ 319] = rx_phy_postflop_0 [ 192];
  assign rx_st_data          [ 320] = rx_phy_postflop_0 [ 193];
  assign rx_st_data          [ 321] = rx_phy_postflop_0 [ 194];
  assign rx_st_data          [ 322] = rx_phy_postflop_0 [ 195];
  assign rx_st_data          [ 323] = rx_phy_postflop_0 [ 196];
  assign rx_st_data          [ 324] = rx_phy_postflop_0 [ 197];
//       DBI                        = rx_phy_postflop_0 [ 198];
//       DBI                        = rx_phy_postflop_0 [ 199];
  assign rx_st_data          [ 325] = rx_phy_postflop_0 [ 200];
  assign rx_st_data          [ 326] = rx_phy_postflop_0 [ 201];
  assign rx_st_data          [ 327] = rx_phy_postflop_0 [ 202];
  assign rx_st_data          [ 328] = rx_phy_postflop_0 [ 203];
  assign rx_st_data          [ 329] = rx_phy_postflop_0 [ 204];
  assign rx_st_data          [ 330] = rx_phy_postflop_0 [ 205];
  assign rx_st_data          [ 331] = rx_phy_postflop_0 [ 206];
  assign rx_st_data          [ 332] = rx_phy_postflop_0 [ 207];
  assign rx_st_data          [ 333] = rx_phy_postflop_0 [ 208];
  assign rx_st_data          [ 334] = rx_phy_postflop_0 [ 209];
  assign rx_st_data          [ 335] = rx_phy_postflop_0 [ 210];
  assign rx_st_data          [ 336] = rx_phy_postflop_0 [ 211];
  assign rx_st_data          [ 337] = rx_phy_postflop_0 [ 212];
  assign rx_st_data          [ 338] = rx_phy_postflop_0 [ 213];
  assign rx_st_data          [ 339] = rx_phy_postflop_0 [ 214];
  assign rx_st_data          [ 340] = rx_phy_postflop_0 [ 215];
  assign rx_st_data          [ 341] = rx_phy_postflop_0 [ 216];
  assign rx_st_data          [ 342] = rx_phy_postflop_0 [ 217];
  assign rx_st_data          [ 343] = rx_phy_postflop_0 [ 218];
  assign rx_st_data          [ 344] = rx_phy_postflop_0 [ 219];
  assign rx_st_data          [ 345] = rx_phy_postflop_0 [ 220];
  assign rx_st_data          [ 346] = rx_phy_postflop_0 [ 221];
  assign rx_st_data          [ 347] = rx_phy_postflop_0 [ 222];
  assign rx_st_data          [ 348] = rx_phy_postflop_0 [ 223];
  assign rx_st_data          [ 349] = rx_phy_postflop_0 [ 224];
  assign rx_st_data          [ 350] = rx_phy_postflop_0 [ 225];
  assign rx_st_data          [ 351] = rx_phy_postflop_0 [ 226];
  assign rx_st_data          [ 352] = rx_phy_postflop_0 [ 227];
  assign rx_st_data          [ 353] = rx_phy_postflop_0 [ 228];
  assign rx_st_data          [ 354] = rx_phy_postflop_0 [ 229];
  assign rx_st_data          [ 355] = rx_phy_postflop_0 [ 230];
  assign rx_st_data          [ 356] = rx_phy_postflop_0 [ 231];
  assign rx_st_data          [ 357] = rx_phy_postflop_0 [ 232];
  assign rx_st_data          [ 358] = rx_phy_postflop_0 [ 233];
  assign rx_st_data          [ 359] = rx_phy_postflop_0 [ 234];
  assign rx_st_data          [ 360] = rx_phy_postflop_0 [ 235];
  assign rx_st_data          [ 361] = rx_phy_postflop_0 [ 236];
  assign rx_st_data          [ 362] = rx_phy_postflop_0 [ 237];
//       DBI                        = rx_phy_postflop_0 [ 238];
//       DBI                        = rx_phy_postflop_0 [ 239];
//       MARKER                     = rx_phy_postflop_1 [ 160]
//       STROBE                     = rx_phy_postflop_1 [ 161]
  assign rx_st_data          [ 363] = rx_phy_postflop_1 [ 162];
  assign rx_st_data          [ 364] = rx_phy_postflop_1 [ 163];
  assign rx_st_data          [ 365] = rx_phy_postflop_1 [ 164];
  assign rx_st_data          [ 366] = rx_phy_postflop_1 [ 165];
  assign rx_st_data          [ 367] = rx_phy_postflop_1 [ 166];
  assign rx_st_data          [ 368] = rx_phy_postflop_1 [ 167];
  assign rx_st_data          [ 369] = rx_phy_postflop_1 [ 168];
  assign rx_st_data          [ 370] = rx_phy_postflop_1 [ 169];
  assign rx_st_data          [ 371] = rx_phy_postflop_1 [ 170];
  assign rx_st_data          [ 372] = rx_phy_postflop_1 [ 171];
  assign rx_st_data          [ 373] = rx_phy_postflop_1 [ 172];
  assign rx_st_data          [ 374] = rx_phy_postflop_1 [ 173];
  assign rx_st_data          [ 375] = rx_phy_postflop_1 [ 174];
  assign rx_st_data          [ 376] = rx_phy_postflop_1 [ 175];
  assign rx_st_data          [ 377] = rx_phy_postflop_1 [ 176];
  assign rx_st_data          [ 378] = rx_phy_postflop_1 [ 177];
  assign rx_st_data          [ 379] = rx_phy_postflop_1 [ 178];
  assign rx_st_data          [ 380] = rx_phy_postflop_1 [ 179];
  assign rx_st_data          [ 381] = rx_phy_postflop_1 [ 180];
  assign rx_st_data          [ 382] = rx_phy_postflop_1 [ 181];
  assign rx_st_data          [ 383] = rx_phy_postflop_1 [ 182];
  assign rx_st_data          [ 384] = rx_phy_postflop_1 [ 183];
  assign rx_st_data          [ 385] = rx_phy_postflop_1 [ 184];
  assign rx_st_data          [ 386] = rx_phy_postflop_1 [ 185];
  assign rx_st_data          [ 387] = rx_phy_postflop_1 [ 186];
  assign rx_st_data          [ 388] = rx_phy_postflop_1 [ 187];
  assign rx_st_data          [ 389] = rx_phy_postflop_1 [ 188];
  assign rx_st_data          [ 390] = rx_phy_postflop_1 [ 189];
  assign rx_st_data          [ 391] = rx_phy_postflop_1 [ 190];
  assign rx_st_data          [ 392] = rx_phy_postflop_1 [ 191];
  assign rx_st_data          [ 393] = rx_phy_postflop_1 [ 192];
  assign rx_st_data          [ 394] = rx_phy_postflop_1 [ 193];
  assign rx_st_data          [ 395] = rx_phy_postflop_1 [ 194];
  assign rx_st_data          [ 396] = rx_phy_postflop_1 [ 195];
  assign rx_st_data          [ 397] = rx_phy_postflop_1 [ 196];
  assign rx_st_data          [ 398] = rx_phy_postflop_1 [ 197];
//       DBI                        = rx_phy_postflop_1 [ 198];
//       DBI                        = rx_phy_postflop_1 [ 199];
  assign rx_st_data          [ 399] = rx_phy_postflop_1 [ 200];
  assign rx_st_data          [ 400] = rx_phy_postflop_1 [ 201];
  assign rx_st_data          [ 401] = rx_phy_postflop_1 [ 202];
  assign rx_st_data          [ 402] = rx_phy_postflop_1 [ 203];
  assign rx_st_data          [ 403] = rx_phy_postflop_1 [ 204];
  assign rx_st_data          [ 404] = rx_phy_postflop_1 [ 205];
  assign rx_st_data          [ 405] = rx_phy_postflop_1 [ 206];
  assign rx_st_data          [ 406] = rx_phy_postflop_1 [ 207];
  assign rx_st_data          [ 407] = rx_phy_postflop_1 [ 208];
  assign rx_st_data          [ 408] = rx_phy_postflop_1 [ 209];
  assign rx_st_data          [ 409] = rx_phy_postflop_1 [ 210];
  assign rx_st_data          [ 410] = rx_phy_postflop_1 [ 211];
  assign rx_st_data          [ 411] = rx_phy_postflop_1 [ 212];
  assign rx_st_data          [ 412] = rx_phy_postflop_1 [ 213];
  assign rx_st_data          [ 413] = rx_phy_postflop_1 [ 214];
  assign rx_st_data          [ 414] = rx_phy_postflop_1 [ 215];
  assign rx_st_data          [ 415] = rx_phy_postflop_1 [ 216];
  assign rx_st_data          [ 416] = rx_phy_postflop_1 [ 217];
  assign rx_st_data          [ 417] = rx_phy_postflop_1 [ 218];
  assign rx_st_data          [ 418] = rx_phy_postflop_1 [ 219];
  assign rx_st_data          [ 419] = rx_phy_postflop_1 [ 220];
  assign rx_st_data          [ 420] = rx_phy_postflop_1 [ 221];
  assign rx_st_data          [ 421] = rx_phy_postflop_1 [ 222];
  assign rx_st_data          [ 422] = rx_phy_postflop_1 [ 223];
  assign rx_st_data          [ 423] = rx_phy_postflop_1 [ 224];
  assign rx_st_data          [ 424] = rx_phy_postflop_1 [ 225];
  assign rx_st_data          [ 425] = rx_phy_postflop_1 [ 226];
  assign rx_st_data          [ 426] = rx_phy_postflop_1 [ 227];
  assign rx_st_data          [ 427] = rx_phy_postflop_1 [ 228];
  assign rx_st_data          [ 428] = rx_phy_postflop_1 [ 229];
  assign rx_st_data          [ 429] = rx_phy_postflop_1 [ 230];
  assign rx_st_data          [ 430] = rx_phy_postflop_1 [ 231];
  assign rx_st_data          [ 431] = rx_phy_postflop_1 [ 232];
  assign rx_st_data          [ 432] = rx_phy_postflop_1 [ 233];
  assign rx_st_data          [ 433] = rx_phy_postflop_1 [ 234];
  assign rx_st_data          [ 434] = rx_phy_postflop_1 [ 235];
//       nc                         = rx_phy_postflop_1 [ 236];
//       nc                         = rx_phy_postflop_1 [ 237];
//       DBI                        = rx_phy_postflop_1 [ 238];
//       DBI                        = rx_phy_postflop_1 [ 239];
//       MARKER                     = rx_phy_postflop_0 [ 240]
//       STROBE                     = rx_phy_postflop_0 [ 241]
  assign rx_st_pushbit_r3           = rx_phy_postflop_0 [ 242];
  assign rx_st_data          [ 435] = rx_phy_postflop_0 [ 243];
  assign rx_st_data          [ 436] = rx_phy_postflop_0 [ 244];
  assign rx_st_data          [ 437] = rx_phy_postflop_0 [ 245];
  assign rx_st_data          [ 438] = rx_phy_postflop_0 [ 246];
  assign rx_st_data          [ 439] = rx_phy_postflop_0 [ 247];
  assign rx_st_data          [ 440] = rx_phy_postflop_0 [ 248];
  assign rx_st_data          [ 441] = rx_phy_postflop_0 [ 249];
  assign rx_st_data          [ 442] = rx_phy_postflop_0 [ 250];
  assign rx_st_data          [ 443] = rx_phy_postflop_0 [ 251];
  assign rx_st_data          [ 444] = rx_phy_postflop_0 [ 252];
  assign rx_st_data          [ 445] = rx_phy_postflop_0 [ 253];
  assign rx_st_data          [ 446] = rx_phy_postflop_0 [ 254];
  assign rx_st_data          [ 447] = rx_phy_postflop_0 [ 255];
  assign rx_st_data          [ 448] = rx_phy_postflop_0 [ 256];
  assign rx_st_data          [ 449] = rx_phy_postflop_0 [ 257];
  assign rx_st_data          [ 450] = rx_phy_postflop_0 [ 258];
  assign rx_st_data          [ 451] = rx_phy_postflop_0 [ 259];
  assign rx_st_data          [ 452] = rx_phy_postflop_0 [ 260];
  assign rx_st_data          [ 453] = rx_phy_postflop_0 [ 261];
  assign rx_st_data          [ 454] = rx_phy_postflop_0 [ 262];
  assign rx_st_data          [ 455] = rx_phy_postflop_0 [ 263];
  assign rx_st_data          [ 456] = rx_phy_postflop_0 [ 264];
  assign rx_st_data          [ 457] = rx_phy_postflop_0 [ 265];
  assign rx_st_data          [ 458] = rx_phy_postflop_0 [ 266];
  assign rx_st_data          [ 459] = rx_phy_postflop_0 [ 267];
  assign rx_st_data          [ 460] = rx_phy_postflop_0 [ 268];
  assign rx_st_data          [ 461] = rx_phy_postflop_0 [ 269];
  assign rx_st_data          [ 462] = rx_phy_postflop_0 [ 270];
  assign rx_st_data          [ 463] = rx_phy_postflop_0 [ 271];
  assign rx_st_data          [ 464] = rx_phy_postflop_0 [ 272];
  assign rx_st_data          [ 465] = rx_phy_postflop_0 [ 273];
  assign rx_st_data          [ 466] = rx_phy_postflop_0 [ 274];
  assign rx_st_data          [ 467] = rx_phy_postflop_0 [ 275];
  assign rx_st_data          [ 468] = rx_phy_postflop_0 [ 276];
  assign rx_st_data          [ 469] = rx_phy_postflop_0 [ 277];
//       DBI                        = rx_phy_postflop_0 [ 278];
//       DBI                        = rx_phy_postflop_0 [ 279];
  assign rx_st_data          [ 470] = rx_phy_postflop_0 [ 280];
  assign rx_st_data          [ 471] = rx_phy_postflop_0 [ 281];
  assign rx_st_data          [ 472] = rx_phy_postflop_0 [ 282];
  assign rx_st_data          [ 473] = rx_phy_postflop_0 [ 283];
  assign rx_st_data          [ 474] = rx_phy_postflop_0 [ 284];
  assign rx_st_data          [ 475] = rx_phy_postflop_0 [ 285];
  assign rx_st_data          [ 476] = rx_phy_postflop_0 [ 286];
  assign rx_st_data          [ 477] = rx_phy_postflop_0 [ 287];
  assign rx_st_data          [ 478] = rx_phy_postflop_0 [ 288];
  assign rx_st_data          [ 479] = rx_phy_postflop_0 [ 289];
  assign rx_st_data          [ 480] = rx_phy_postflop_0 [ 290];
  assign rx_st_data          [ 481] = rx_phy_postflop_0 [ 291];
  assign rx_st_data          [ 482] = rx_phy_postflop_0 [ 292];
  assign rx_st_data          [ 483] = rx_phy_postflop_0 [ 293];
  assign rx_st_data          [ 484] = rx_phy_postflop_0 [ 294];
  assign rx_st_data          [ 485] = rx_phy_postflop_0 [ 295];
  assign rx_st_data          [ 486] = rx_phy_postflop_0 [ 296];
  assign rx_st_data          [ 487] = rx_phy_postflop_0 [ 297];
  assign rx_st_data          [ 488] = rx_phy_postflop_0 [ 298];
  assign rx_st_data          [ 489] = rx_phy_postflop_0 [ 299];
  assign rx_st_data          [ 490] = rx_phy_postflop_0 [ 300];
  assign rx_st_data          [ 491] = rx_phy_postflop_0 [ 301];
  assign rx_st_data          [ 492] = rx_phy_postflop_0 [ 302];
  assign rx_st_data          [ 493] = rx_phy_postflop_0 [ 303];
  assign rx_st_data          [ 494] = rx_phy_postflop_0 [ 304];
  assign rx_st_data          [ 495] = rx_phy_postflop_0 [ 305];
  assign rx_st_data          [ 496] = rx_phy_postflop_0 [ 306];
  assign rx_st_data          [ 497] = rx_phy_postflop_0 [ 307];
  assign rx_st_data          [ 498] = rx_phy_postflop_0 [ 308];
  assign rx_st_data          [ 499] = rx_phy_postflop_0 [ 309];
  assign rx_st_data          [ 500] = rx_phy_postflop_0 [ 310];
  assign rx_st_data          [ 501] = rx_phy_postflop_0 [ 311];
  assign rx_st_data          [ 502] = rx_phy_postflop_0 [ 312];
  assign rx_st_data          [ 503] = rx_phy_postflop_0 [ 313];
  assign rx_st_data          [ 504] = rx_phy_postflop_0 [ 314];
  assign rx_st_data          [ 505] = rx_phy_postflop_0 [ 315];
  assign rx_st_data          [ 506] = rx_phy_postflop_0 [ 316];
  assign rx_st_data          [ 507] = rx_phy_postflop_0 [ 317];
//       DBI                        = rx_phy_postflop_0 [ 318];
//       DBI                        = rx_phy_postflop_0 [ 319];
//       MARKER                     = rx_phy_postflop_1 [ 240]
//       STROBE                     = rx_phy_postflop_1 [ 241]
  assign rx_st_data          [ 508] = rx_phy_postflop_1 [ 242];
  assign rx_st_data          [ 509] = rx_phy_postflop_1 [ 243];
  assign rx_st_data          [ 510] = rx_phy_postflop_1 [ 244];
  assign rx_st_data          [ 511] = rx_phy_postflop_1 [ 245];
  assign rx_st_data          [ 512] = rx_phy_postflop_1 [ 246];
  assign rx_st_data          [ 513] = rx_phy_postflop_1 [ 247];
  assign rx_st_data          [ 514] = rx_phy_postflop_1 [ 248];
  assign rx_st_data          [ 515] = rx_phy_postflop_1 [ 249];
  assign rx_st_data          [ 516] = rx_phy_postflop_1 [ 250];
  assign rx_st_data          [ 517] = rx_phy_postflop_1 [ 251];
  assign rx_st_data          [ 518] = rx_phy_postflop_1 [ 252];
  assign rx_st_data          [ 519] = rx_phy_postflop_1 [ 253];
  assign rx_st_data          [ 520] = rx_phy_postflop_1 [ 254];
  assign rx_st_data          [ 521] = rx_phy_postflop_1 [ 255];
  assign rx_st_data          [ 522] = rx_phy_postflop_1 [ 256];
  assign rx_st_data          [ 523] = rx_phy_postflop_1 [ 257];
  assign rx_st_data          [ 524] = rx_phy_postflop_1 [ 258];
  assign rx_st_data          [ 525] = rx_phy_postflop_1 [ 259];
  assign rx_st_data          [ 526] = rx_phy_postflop_1 [ 260];
  assign rx_st_data          [ 527] = rx_phy_postflop_1 [ 261];
  assign rx_st_data          [ 528] = rx_phy_postflop_1 [ 262];
  assign rx_st_data          [ 529] = rx_phy_postflop_1 [ 263];
  assign rx_st_data          [ 530] = rx_phy_postflop_1 [ 264];
  assign rx_st_data          [ 531] = rx_phy_postflop_1 [ 265];
  assign rx_st_data          [ 532] = rx_phy_postflop_1 [ 266];
  assign rx_st_data          [ 533] = rx_phy_postflop_1 [ 267];
  assign rx_st_data          [ 534] = rx_phy_postflop_1 [ 268];
  assign rx_st_data          [ 535] = rx_phy_postflop_1 [ 269];
  assign rx_st_data          [ 536] = rx_phy_postflop_1 [ 270];
  assign rx_st_data          [ 537] = rx_phy_postflop_1 [ 271];
  assign rx_st_data          [ 538] = rx_phy_postflop_1 [ 272];
  assign rx_st_data          [ 539] = rx_phy_postflop_1 [ 273];
  assign rx_st_data          [ 540] = rx_phy_postflop_1 [ 274];
  assign rx_st_data          [ 541] = rx_phy_postflop_1 [ 275];
  assign rx_st_data          [ 542] = rx_phy_postflop_1 [ 276];
  assign rx_st_data          [ 543] = rx_phy_postflop_1 [ 277];
//       DBI                        = rx_phy_postflop_1 [ 278];
//       DBI                        = rx_phy_postflop_1 [ 279];
  assign rx_st_data          [ 544] = rx_phy_postflop_1 [ 280];
  assign rx_st_data          [ 545] = rx_phy_postflop_1 [ 281];
  assign rx_st_data          [ 546] = rx_phy_postflop_1 [ 282];
  assign rx_st_data          [ 547] = rx_phy_postflop_1 [ 283];
  assign rx_st_data          [ 548] = rx_phy_postflop_1 [ 284];
  assign rx_st_data          [ 549] = rx_phy_postflop_1 [ 285];
  assign rx_st_data          [ 550] = rx_phy_postflop_1 [ 286];
  assign rx_st_data          [ 551] = rx_phy_postflop_1 [ 287];
  assign rx_st_data          [ 552] = rx_phy_postflop_1 [ 288];
  assign rx_st_data          [ 553] = rx_phy_postflop_1 [ 289];
  assign rx_st_data          [ 554] = rx_phy_postflop_1 [ 290];
  assign rx_st_data          [ 555] = rx_phy_postflop_1 [ 291];
  assign rx_st_data          [ 556] = rx_phy_postflop_1 [ 292];
  assign rx_st_data          [ 557] = rx_phy_postflop_1 [ 293];
  assign rx_st_data          [ 558] = rx_phy_postflop_1 [ 294];
  assign rx_st_data          [ 559] = rx_phy_postflop_1 [ 295];
  assign rx_st_data          [ 560] = rx_phy_postflop_1 [ 296];
  assign rx_st_data          [ 561] = rx_phy_postflop_1 [ 297];
  assign rx_st_data          [ 562] = rx_phy_postflop_1 [ 298];
  assign rx_st_data          [ 563] = rx_phy_postflop_1 [ 299];
  assign rx_st_data          [ 564] = rx_phy_postflop_1 [ 300];
  assign rx_st_data          [ 565] = rx_phy_postflop_1 [ 301];
  assign rx_st_data          [ 566] = rx_phy_postflop_1 [ 302];
  assign rx_st_data          [ 567] = rx_phy_postflop_1 [ 303];
  assign rx_st_data          [ 568] = rx_phy_postflop_1 [ 304];
  assign rx_st_data          [ 569] = rx_phy_postflop_1 [ 305];
  assign rx_st_data          [ 570] = rx_phy_postflop_1 [ 306];
  assign rx_st_data          [ 571] = rx_phy_postflop_1 [ 307];
  assign rx_st_data          [ 572] = rx_phy_postflop_1 [ 308];
  assign rx_st_data          [ 573] = rx_phy_postflop_1 [ 309];
  assign rx_st_data          [ 574] = rx_phy_postflop_1 [ 310];
  assign rx_st_data          [ 575] = rx_phy_postflop_1 [ 311];
  assign rx_st_data          [ 576] = rx_phy_postflop_1 [ 312];
  assign rx_st_data          [ 577] = rx_phy_postflop_1 [ 313];
  assign rx_st_data          [ 578] = rx_phy_postflop_1 [ 314];
  assign rx_st_data          [ 579] = rx_phy_postflop_1 [ 315];
//       nc                         = rx_phy_postflop_1 [ 316];
//       nc                         = rx_phy_postflop_1 [ 317];
//       DBI                        = rx_phy_postflop_1 [ 318];
//       DBI                        = rx_phy_postflop_1 [ 319];
  assign rx_st_data          [ 580] = rx_st_pushbit_r0;
  assign rx_st_data          [ 581] = rx_st_pushbit_r1;
  assign rx_st_data          [ 582] = rx_st_pushbit_r2;
  assign rx_st_data          [ 583] = rx_st_pushbit_r3;

// RX Section
//////////////////////////////////////////////////////////////////


endmodule
