////////////////////////////////////////////////////////////
// Proprietary Information of Eximius Design
//
//        (C) Copyright 2021 Eximius Design
//                All Rights Reserved
//
// This entire notice must be reproduced on all copies of this file
// and copies of this file may only be made by a person if such person is
// permitted to do so under the terms of a subsisting license agreement
// from Eximius Design
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
////////////////////////////////////////////////////////////

module axi_st_d128_asym_quarter_master_concat  (

// Data from Logic Links
  input  logic [ 579:   0]   tx_st_data          ,
  output logic               tx_st_pop_ovrd      ,
  input  logic               tx_st_pushbit       ,
  output logic [   3:   0]   rx_st_credit        ,

// PHY Interconnect
  output logic [ 319:   0]   tx_phy0             ,
  input  logic [ 319:   0]   rx_phy0             ,
  output logic [ 319:   0]   tx_phy1             ,
  input  logic [ 319:   0]   rx_phy1             ,

  input  logic               clk_wr              ,
  input  logic               clk_rd              ,
  input  logic               rst_wr_n            ,
  input  logic               rst_rd_n            ,

  input  logic               m_gen2_mode         ,
  input  logic               tx_online           ,

  input  logic               tx_stb_userbit      ,
  input  logic [   3:   0]   tx_mrk_userbit      

);

// No TX Packetization, so tie off packetization signals
  assign tx_st_pop_ovrd                     = 1'b0                               ;

// No RX Packetization, so tie off packetization signals

//////////////////////////////////////////////////////////////////
// TX Section

//   TX_CH_WIDTH           = 320; // Gen2Only running at Quarter Rate
//   TX_DATA_WIDTH         = 296; // Usable Data per Channel
//   TX_PERSISTENT_STROBE  = 1'b1;
//   TX_PERSISTENT_MARKER  = 1'b1;
//   TX_STROBE_GEN2_LOC    = 'd1;
//   TX_MARKER_GEN2_LOC    = 'd0;
//   TX_STROBE_GEN1_LOC    = 'd38;
//   TX_MARKER_GEN1_LOC    = 'd39;
//   TX_ENABLE_STROBE      = 1'b1;
//   TX_ENABLE_MARKER      = 1'b1;
//   TX_DBI_PRESENT        = 1'b1;
//   TX_REG_PHY            = 1'b0;

  localparam TX_REG_PHY    = 1'b0;  // If set, this enables boundary FF for timing reasons

  logic [ 319:   0]                              tx_phy_preflop_0              ;
  logic [ 319:   0]                              tx_phy_preflop_1              ;
  logic [ 319:   0]                              tx_phy_flop_0_reg             ;
  logic [ 319:   0]                              tx_phy_flop_1_reg             ;

  always_ff @(posedge clk_wr or negedge rst_wr_n)
  if (~rst_wr_n)
  begin
    tx_phy_flop_0_reg                       <= 320'b0                                  ;
    tx_phy_flop_1_reg                       <= 320'b0                                  ;
  end
  else
  begin
    tx_phy_flop_0_reg                       <= tx_phy_preflop_0                        ;
    tx_phy_flop_1_reg                       <= tx_phy_preflop_1                        ;
  end

  assign tx_phy0                            = TX_REG_PHY ? tx_phy_flop_0_reg : tx_phy_preflop_0               ;
  assign tx_phy1                            = TX_REG_PHY ? tx_phy_flop_1_reg : tx_phy_preflop_1               ;

  logic                                          tx_st_pushbit_r0              ;
  logic                                          tx_st_pushbit_r1              ;
  logic                                          tx_st_pushbit_r2              ;
  logic                                          tx_st_pushbit_r3              ;

  assign tx_st_pushbit_r0                   = tx_st_pushbit                      ;
  assign tx_st_pushbit_r1                   = tx_st_pushbit                      ;
  assign tx_st_pushbit_r2                   = tx_st_pushbit                      ;
  assign tx_st_pushbit_r3                   = tx_st_pushbit                      ;

  assign tx_phy_preflop_0 [   0] = tx_mrk_userbit[0]          ; // MARKER
  assign tx_phy_preflop_0 [   1] = tx_stb_userbit             ; // STROBE
  assign tx_phy_preflop_0 [   2] = tx_st_pushbit_r0           ;
  assign tx_phy_preflop_0 [   3] = tx_st_data          [   0] ;
  assign tx_phy_preflop_0 [   4] = tx_st_data          [   1] ;
  assign tx_phy_preflop_0 [   5] = tx_st_data          [   2] ;
  assign tx_phy_preflop_0 [   6] = tx_st_data          [   3] ;
  assign tx_phy_preflop_0 [   7] = tx_st_data          [   4] ;
  assign tx_phy_preflop_0 [   8] = tx_st_data          [   5] ;
  assign tx_phy_preflop_0 [   9] = tx_st_data          [   6] ;
  assign tx_phy_preflop_0 [  10] = tx_st_data          [   7] ;
  assign tx_phy_preflop_0 [  11] = tx_st_data          [   8] ;
  assign tx_phy_preflop_0 [  12] = tx_st_data          [   9] ;
  assign tx_phy_preflop_0 [  13] = tx_st_data          [  10] ;
  assign tx_phy_preflop_0 [  14] = tx_st_data          [  11] ;
  assign tx_phy_preflop_0 [  15] = tx_st_data          [  12] ;
  assign tx_phy_preflop_0 [  16] = tx_st_data          [  13] ;
  assign tx_phy_preflop_0 [  17] = tx_st_data          [  14] ;
  assign tx_phy_preflop_0 [  18] = tx_st_data          [  15] ;
  assign tx_phy_preflop_0 [  19] = tx_st_data          [  16] ;
  assign tx_phy_preflop_0 [  20] = tx_st_data          [  17] ;
  assign tx_phy_preflop_0 [  21] = tx_st_data          [  18] ;
  assign tx_phy_preflop_0 [  22] = tx_st_data          [  19] ;
  assign tx_phy_preflop_0 [  23] = tx_st_data          [  20] ;
  assign tx_phy_preflop_0 [  24] = tx_st_data          [  21] ;
  assign tx_phy_preflop_0 [  25] = tx_st_data          [  22] ;
  assign tx_phy_preflop_0 [  26] = tx_st_data          [  23] ;
  assign tx_phy_preflop_0 [  27] = tx_st_data          [  24] ;
  assign tx_phy_preflop_0 [  28] = tx_st_data          [  25] ;
  assign tx_phy_preflop_0 [  29] = tx_st_data          [  26] ;
  assign tx_phy_preflop_0 [  30] = tx_st_data          [  27] ;
  assign tx_phy_preflop_0 [  31] = tx_st_data          [  28] ;
  assign tx_phy_preflop_0 [  32] = tx_st_data          [  29] ;
  assign tx_phy_preflop_0 [  33] = tx_st_data          [  30] ;
  assign tx_phy_preflop_0 [  34] = tx_st_data          [  31] ;
  assign tx_phy_preflop_0 [  35] = tx_st_data          [  32] ;
  assign tx_phy_preflop_0 [  36] = tx_st_data          [  33] ;
  assign tx_phy_preflop_0 [  37] = tx_st_data          [  34] ;
  assign tx_phy_preflop_0 [  38] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [  39] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [  40] = tx_st_data          [  35] ;
  assign tx_phy_preflop_0 [  41] = tx_st_data          [  36] ;
  assign tx_phy_preflop_0 [  42] = tx_st_data          [  37] ;
  assign tx_phy_preflop_0 [  43] = tx_st_data          [  38] ;
  assign tx_phy_preflop_0 [  44] = tx_st_data          [  39] ;
  assign tx_phy_preflop_0 [  45] = tx_st_data          [  40] ;
  assign tx_phy_preflop_0 [  46] = tx_st_data          [  41] ;
  assign tx_phy_preflop_0 [  47] = tx_st_data          [  42] ;
  assign tx_phy_preflop_0 [  48] = tx_st_data          [  43] ;
  assign tx_phy_preflop_0 [  49] = tx_st_data          [  44] ;
  assign tx_phy_preflop_0 [  50] = tx_st_data          [  45] ;
  assign tx_phy_preflop_0 [  51] = tx_st_data          [  46] ;
  assign tx_phy_preflop_0 [  52] = tx_st_data          [  47] ;
  assign tx_phy_preflop_0 [  53] = tx_st_data          [  48] ;
  assign tx_phy_preflop_0 [  54] = tx_st_data          [  49] ;
  assign tx_phy_preflop_0 [  55] = tx_st_data          [  50] ;
  assign tx_phy_preflop_0 [  56] = tx_st_data          [  51] ;
  assign tx_phy_preflop_0 [  57] = tx_st_data          [  52] ;
  assign tx_phy_preflop_0 [  58] = tx_st_data          [  53] ;
  assign tx_phy_preflop_0 [  59] = tx_st_data          [  54] ;
  assign tx_phy_preflop_0 [  60] = tx_st_data          [  55] ;
  assign tx_phy_preflop_0 [  61] = tx_st_data          [  56] ;
  assign tx_phy_preflop_0 [  62] = tx_st_data          [  57] ;
  assign tx_phy_preflop_0 [  63] = tx_st_data          [  58] ;
  assign tx_phy_preflop_0 [  64] = tx_st_data          [  59] ;
  assign tx_phy_preflop_0 [  65] = tx_st_data          [  60] ;
  assign tx_phy_preflop_0 [  66] = tx_st_data          [  61] ;
  assign tx_phy_preflop_0 [  67] = tx_st_data          [  62] ;
  assign tx_phy_preflop_0 [  68] = tx_st_data          [  63] ;
  assign tx_phy_preflop_0 [  69] = tx_st_data          [  64] ;
  assign tx_phy_preflop_0 [  70] = tx_st_data          [  65] ;
  assign tx_phy_preflop_0 [  71] = tx_st_data          [  66] ;
  assign tx_phy_preflop_0 [  72] = tx_st_data          [  67] ;
  assign tx_phy_preflop_0 [  73] = tx_st_data          [  68] ;
  assign tx_phy_preflop_0 [  74] = tx_st_data          [  69] ;
  assign tx_phy_preflop_0 [  75] = tx_st_data          [  70] ;
  assign tx_phy_preflop_0 [  76] = tx_st_data          [  71] ;
  assign tx_phy_preflop_0 [  77] = tx_st_data          [  72] ;
  assign tx_phy_preflop_0 [  78] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [  79] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [   0] = tx_mrk_userbit[0]          ; // MARKER
  assign tx_phy_preflop_1 [   1] = tx_stb_userbit             ; // STROBE
  assign tx_phy_preflop_1 [   2] = tx_st_data          [  73] ;
  assign tx_phy_preflop_1 [   3] = tx_st_data          [  74] ;
  assign tx_phy_preflop_1 [   4] = tx_st_data          [  75] ;
  assign tx_phy_preflop_1 [   5] = tx_st_data          [  76] ;
  assign tx_phy_preflop_1 [   6] = tx_st_data          [  77] ;
  assign tx_phy_preflop_1 [   7] = tx_st_data          [  78] ;
  assign tx_phy_preflop_1 [   8] = tx_st_data          [  79] ;
  assign tx_phy_preflop_1 [   9] = tx_st_data          [  80] ;
  assign tx_phy_preflop_1 [  10] = tx_st_data          [  81] ;
  assign tx_phy_preflop_1 [  11] = tx_st_data          [  82] ;
  assign tx_phy_preflop_1 [  12] = tx_st_data          [  83] ;
  assign tx_phy_preflop_1 [  13] = tx_st_data          [  84] ;
  assign tx_phy_preflop_1 [  14] = tx_st_data          [  85] ;
  assign tx_phy_preflop_1 [  15] = tx_st_data          [  86] ;
  assign tx_phy_preflop_1 [  16] = tx_st_data          [  87] ;
  assign tx_phy_preflop_1 [  17] = tx_st_data          [  88] ;
  assign tx_phy_preflop_1 [  18] = tx_st_data          [  89] ;
  assign tx_phy_preflop_1 [  19] = tx_st_data          [  90] ;
  assign tx_phy_preflop_1 [  20] = tx_st_data          [  91] ;
  assign tx_phy_preflop_1 [  21] = tx_st_data          [  92] ;
  assign tx_phy_preflop_1 [  22] = tx_st_data          [  93] ;
  assign tx_phy_preflop_1 [  23] = tx_st_data          [  94] ;
  assign tx_phy_preflop_1 [  24] = tx_st_data          [  95] ;
  assign tx_phy_preflop_1 [  25] = tx_st_data          [  96] ;
  assign tx_phy_preflop_1 [  26] = tx_st_data          [  97] ;
  assign tx_phy_preflop_1 [  27] = tx_st_data          [  98] ;
  assign tx_phy_preflop_1 [  28] = tx_st_data          [  99] ;
  assign tx_phy_preflop_1 [  29] = tx_st_data          [ 100] ;
  assign tx_phy_preflop_1 [  30] = tx_st_data          [ 101] ;
  assign tx_phy_preflop_1 [  31] = tx_st_data          [ 102] ;
  assign tx_phy_preflop_1 [  32] = tx_st_data          [ 103] ;
  assign tx_phy_preflop_1 [  33] = tx_st_data          [ 104] ;
  assign tx_phy_preflop_1 [  34] = tx_st_data          [ 105] ;
  assign tx_phy_preflop_1 [  35] = tx_st_data          [ 106] ;
  assign tx_phy_preflop_1 [  36] = tx_st_data          [ 107] ;
  assign tx_phy_preflop_1 [  37] = tx_st_data          [ 108] ;
  assign tx_phy_preflop_1 [  38] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [  39] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [  40] = tx_st_data          [ 109] ;
  assign tx_phy_preflop_1 [  41] = tx_st_data          [ 110] ;
  assign tx_phy_preflop_1 [  42] = tx_st_data          [ 111] ;
  assign tx_phy_preflop_1 [  43] = tx_st_data          [ 112] ;
  assign tx_phy_preflop_1 [  44] = tx_st_data          [ 113] ;
  assign tx_phy_preflop_1 [  45] = tx_st_data          [ 114] ;
  assign tx_phy_preflop_1 [  46] = tx_st_data          [ 115] ;
  assign tx_phy_preflop_1 [  47] = tx_st_data          [ 116] ;
  assign tx_phy_preflop_1 [  48] = tx_st_data          [ 117] ;
  assign tx_phy_preflop_1 [  49] = tx_st_data          [ 118] ;
  assign tx_phy_preflop_1 [  50] = tx_st_data          [ 119] ;
  assign tx_phy_preflop_1 [  51] = tx_st_data          [ 120] ;
  assign tx_phy_preflop_1 [  52] = tx_st_data          [ 121] ;
  assign tx_phy_preflop_1 [  53] = tx_st_data          [ 122] ;
  assign tx_phy_preflop_1 [  54] = tx_st_data          [ 123] ;
  assign tx_phy_preflop_1 [  55] = tx_st_data          [ 124] ;
  assign tx_phy_preflop_1 [  56] = tx_st_data          [ 125] ;
  assign tx_phy_preflop_1 [  57] = tx_st_data          [ 126] ;
  assign tx_phy_preflop_1 [  58] = tx_st_data          [ 127] ;
  assign tx_phy_preflop_1 [  59] = tx_st_data          [ 128] ;
  assign tx_phy_preflop_1 [  60] = tx_st_data          [ 129] ;
  assign tx_phy_preflop_1 [  61] = tx_st_data          [ 130] ;
  assign tx_phy_preflop_1 [  62] = tx_st_data          [ 131] ;
  assign tx_phy_preflop_1 [  63] = tx_st_data          [ 132] ;
  assign tx_phy_preflop_1 [  64] = tx_st_data          [ 133] ;
  assign tx_phy_preflop_1 [  65] = tx_st_data          [ 134] ;
  assign tx_phy_preflop_1 [  66] = tx_st_data          [ 135] ;
  assign tx_phy_preflop_1 [  67] = tx_st_data          [ 136] ;
  assign tx_phy_preflop_1 [  68] = tx_st_data          [ 137] ;
  assign tx_phy_preflop_1 [  69] = tx_st_data          [ 138] ;
  assign tx_phy_preflop_1 [  70] = tx_st_data          [ 139] ;
  assign tx_phy_preflop_1 [  71] = tx_st_data          [ 140] ;
  assign tx_phy_preflop_1 [  72] = tx_st_data          [ 141] ;
  assign tx_phy_preflop_1 [  73] = tx_st_data          [ 142] ;
  assign tx_phy_preflop_1 [  74] = tx_st_data          [ 143] ;
  assign tx_phy_preflop_1 [  75] = tx_st_data          [ 144] ;
  assign tx_phy_preflop_1 [  76] = 1'b0                       ;
  assign tx_phy_preflop_1 [  77] = 1'b0                       ;
  assign tx_phy_preflop_1 [  78] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [  79] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [  80] = tx_mrk_userbit[1]          ; // MARKER
  assign tx_phy_preflop_0 [  81] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_0 [  82] = tx_st_pushbit_r1           ;
  assign tx_phy_preflop_0 [  83] = tx_st_data          [ 145] ;
  assign tx_phy_preflop_0 [  84] = tx_st_data          [ 146] ;
  assign tx_phy_preflop_0 [  85] = tx_st_data          [ 147] ;
  assign tx_phy_preflop_0 [  86] = tx_st_data          [ 148] ;
  assign tx_phy_preflop_0 [  87] = tx_st_data          [ 149] ;
  assign tx_phy_preflop_0 [  88] = tx_st_data          [ 150] ;
  assign tx_phy_preflop_0 [  89] = tx_st_data          [ 151] ;
  assign tx_phy_preflop_0 [  90] = tx_st_data          [ 152] ;
  assign tx_phy_preflop_0 [  91] = tx_st_data          [ 153] ;
  assign tx_phy_preflop_0 [  92] = tx_st_data          [ 154] ;
  assign tx_phy_preflop_0 [  93] = tx_st_data          [ 155] ;
  assign tx_phy_preflop_0 [  94] = tx_st_data          [ 156] ;
  assign tx_phy_preflop_0 [  95] = tx_st_data          [ 157] ;
  assign tx_phy_preflop_0 [  96] = tx_st_data          [ 158] ;
  assign tx_phy_preflop_0 [  97] = tx_st_data          [ 159] ;
  assign tx_phy_preflop_0 [  98] = tx_st_data          [ 160] ;
  assign tx_phy_preflop_0 [  99] = tx_st_data          [ 161] ;
  assign tx_phy_preflop_0 [ 100] = tx_st_data          [ 162] ;
  assign tx_phy_preflop_0 [ 101] = tx_st_data          [ 163] ;
  assign tx_phy_preflop_0 [ 102] = tx_st_data          [ 164] ;
  assign tx_phy_preflop_0 [ 103] = tx_st_data          [ 165] ;
  assign tx_phy_preflop_0 [ 104] = tx_st_data          [ 166] ;
  assign tx_phy_preflop_0 [ 105] = tx_st_data          [ 167] ;
  assign tx_phy_preflop_0 [ 106] = tx_st_data          [ 168] ;
  assign tx_phy_preflop_0 [ 107] = tx_st_data          [ 169] ;
  assign tx_phy_preflop_0 [ 108] = tx_st_data          [ 170] ;
  assign tx_phy_preflop_0 [ 109] = tx_st_data          [ 171] ;
  assign tx_phy_preflop_0 [ 110] = tx_st_data          [ 172] ;
  assign tx_phy_preflop_0 [ 111] = tx_st_data          [ 173] ;
  assign tx_phy_preflop_0 [ 112] = tx_st_data          [ 174] ;
  assign tx_phy_preflop_0 [ 113] = tx_st_data          [ 175] ;
  assign tx_phy_preflop_0 [ 114] = tx_st_data          [ 176] ;
  assign tx_phy_preflop_0 [ 115] = tx_st_data          [ 177] ;
  assign tx_phy_preflop_0 [ 116] = tx_st_data          [ 178] ;
  assign tx_phy_preflop_0 [ 117] = tx_st_data          [ 179] ;
  assign tx_phy_preflop_0 [ 118] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 119] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 120] = tx_st_data          [ 180] ;
  assign tx_phy_preflop_0 [ 121] = tx_st_data          [ 181] ;
  assign tx_phy_preflop_0 [ 122] = tx_st_data          [ 182] ;
  assign tx_phy_preflop_0 [ 123] = tx_st_data          [ 183] ;
  assign tx_phy_preflop_0 [ 124] = tx_st_data          [ 184] ;
  assign tx_phy_preflop_0 [ 125] = tx_st_data          [ 185] ;
  assign tx_phy_preflop_0 [ 126] = tx_st_data          [ 186] ;
  assign tx_phy_preflop_0 [ 127] = tx_st_data          [ 187] ;
  assign tx_phy_preflop_0 [ 128] = tx_st_data          [ 188] ;
  assign tx_phy_preflop_0 [ 129] = tx_st_data          [ 189] ;
  assign tx_phy_preflop_0 [ 130] = tx_st_data          [ 190] ;
  assign tx_phy_preflop_0 [ 131] = tx_st_data          [ 191] ;
  assign tx_phy_preflop_0 [ 132] = tx_st_data          [ 192] ;
  assign tx_phy_preflop_0 [ 133] = tx_st_data          [ 193] ;
  assign tx_phy_preflop_0 [ 134] = tx_st_data          [ 194] ;
  assign tx_phy_preflop_0 [ 135] = tx_st_data          [ 195] ;
  assign tx_phy_preflop_0 [ 136] = tx_st_data          [ 196] ;
  assign tx_phy_preflop_0 [ 137] = tx_st_data          [ 197] ;
  assign tx_phy_preflop_0 [ 138] = tx_st_data          [ 198] ;
  assign tx_phy_preflop_0 [ 139] = tx_st_data          [ 199] ;
  assign tx_phy_preflop_0 [ 140] = tx_st_data          [ 200] ;
  assign tx_phy_preflop_0 [ 141] = tx_st_data          [ 201] ;
  assign tx_phy_preflop_0 [ 142] = tx_st_data          [ 202] ;
  assign tx_phy_preflop_0 [ 143] = tx_st_data          [ 203] ;
  assign tx_phy_preflop_0 [ 144] = tx_st_data          [ 204] ;
  assign tx_phy_preflop_0 [ 145] = tx_st_data          [ 205] ;
  assign tx_phy_preflop_0 [ 146] = tx_st_data          [ 206] ;
  assign tx_phy_preflop_0 [ 147] = tx_st_data          [ 207] ;
  assign tx_phy_preflop_0 [ 148] = tx_st_data          [ 208] ;
  assign tx_phy_preflop_0 [ 149] = tx_st_data          [ 209] ;
  assign tx_phy_preflop_0 [ 150] = tx_st_data          [ 210] ;
  assign tx_phy_preflop_0 [ 151] = tx_st_data          [ 211] ;
  assign tx_phy_preflop_0 [ 152] = tx_st_data          [ 212] ;
  assign tx_phy_preflop_0 [ 153] = tx_st_data          [ 213] ;
  assign tx_phy_preflop_0 [ 154] = tx_st_data          [ 214] ;
  assign tx_phy_preflop_0 [ 155] = tx_st_data          [ 215] ;
  assign tx_phy_preflop_0 [ 156] = tx_st_data          [ 216] ;
  assign tx_phy_preflop_0 [ 157] = tx_st_data          [ 217] ;
  assign tx_phy_preflop_0 [ 158] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 159] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [  80] = tx_mrk_userbit[1]          ; // MARKER
  assign tx_phy_preflop_1 [  81] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_1 [  82] = tx_st_data          [ 218] ;
  assign tx_phy_preflop_1 [  83] = tx_st_data          [ 219] ;
  assign tx_phy_preflop_1 [  84] = tx_st_data          [ 220] ;
  assign tx_phy_preflop_1 [  85] = tx_st_data          [ 221] ;
  assign tx_phy_preflop_1 [  86] = tx_st_data          [ 222] ;
  assign tx_phy_preflop_1 [  87] = tx_st_data          [ 223] ;
  assign tx_phy_preflop_1 [  88] = tx_st_data          [ 224] ;
  assign tx_phy_preflop_1 [  89] = tx_st_data          [ 225] ;
  assign tx_phy_preflop_1 [  90] = tx_st_data          [ 226] ;
  assign tx_phy_preflop_1 [  91] = tx_st_data          [ 227] ;
  assign tx_phy_preflop_1 [  92] = tx_st_data          [ 228] ;
  assign tx_phy_preflop_1 [  93] = tx_st_data          [ 229] ;
  assign tx_phy_preflop_1 [  94] = tx_st_data          [ 230] ;
  assign tx_phy_preflop_1 [  95] = tx_st_data          [ 231] ;
  assign tx_phy_preflop_1 [  96] = tx_st_data          [ 232] ;
  assign tx_phy_preflop_1 [  97] = tx_st_data          [ 233] ;
  assign tx_phy_preflop_1 [  98] = tx_st_data          [ 234] ;
  assign tx_phy_preflop_1 [  99] = tx_st_data          [ 235] ;
  assign tx_phy_preflop_1 [ 100] = tx_st_data          [ 236] ;
  assign tx_phy_preflop_1 [ 101] = tx_st_data          [ 237] ;
  assign tx_phy_preflop_1 [ 102] = tx_st_data          [ 238] ;
  assign tx_phy_preflop_1 [ 103] = tx_st_data          [ 239] ;
  assign tx_phy_preflop_1 [ 104] = tx_st_data          [ 240] ;
  assign tx_phy_preflop_1 [ 105] = tx_st_data          [ 241] ;
  assign tx_phy_preflop_1 [ 106] = tx_st_data          [ 242] ;
  assign tx_phy_preflop_1 [ 107] = tx_st_data          [ 243] ;
  assign tx_phy_preflop_1 [ 108] = tx_st_data          [ 244] ;
  assign tx_phy_preflop_1 [ 109] = tx_st_data          [ 245] ;
  assign tx_phy_preflop_1 [ 110] = tx_st_data          [ 246] ;
  assign tx_phy_preflop_1 [ 111] = tx_st_data          [ 247] ;
  assign tx_phy_preflop_1 [ 112] = tx_st_data          [ 248] ;
  assign tx_phy_preflop_1 [ 113] = tx_st_data          [ 249] ;
  assign tx_phy_preflop_1 [ 114] = tx_st_data          [ 250] ;
  assign tx_phy_preflop_1 [ 115] = tx_st_data          [ 251] ;
  assign tx_phy_preflop_1 [ 116] = tx_st_data          [ 252] ;
  assign tx_phy_preflop_1 [ 117] = tx_st_data          [ 253] ;
  assign tx_phy_preflop_1 [ 118] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 119] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 120] = tx_st_data          [ 254] ;
  assign tx_phy_preflop_1 [ 121] = tx_st_data          [ 255] ;
  assign tx_phy_preflop_1 [ 122] = tx_st_data          [ 256] ;
  assign tx_phy_preflop_1 [ 123] = tx_st_data          [ 257] ;
  assign tx_phy_preflop_1 [ 124] = tx_st_data          [ 258] ;
  assign tx_phy_preflop_1 [ 125] = tx_st_data          [ 259] ;
  assign tx_phy_preflop_1 [ 126] = tx_st_data          [ 260] ;
  assign tx_phy_preflop_1 [ 127] = tx_st_data          [ 261] ;
  assign tx_phy_preflop_1 [ 128] = tx_st_data          [ 262] ;
  assign tx_phy_preflop_1 [ 129] = tx_st_data          [ 263] ;
  assign tx_phy_preflop_1 [ 130] = tx_st_data          [ 264] ;
  assign tx_phy_preflop_1 [ 131] = tx_st_data          [ 265] ;
  assign tx_phy_preflop_1 [ 132] = tx_st_data          [ 266] ;
  assign tx_phy_preflop_1 [ 133] = tx_st_data          [ 267] ;
  assign tx_phy_preflop_1 [ 134] = tx_st_data          [ 268] ;
  assign tx_phy_preflop_1 [ 135] = tx_st_data          [ 269] ;
  assign tx_phy_preflop_1 [ 136] = tx_st_data          [ 270] ;
  assign tx_phy_preflop_1 [ 137] = tx_st_data          [ 271] ;
  assign tx_phy_preflop_1 [ 138] = tx_st_data          [ 272] ;
  assign tx_phy_preflop_1 [ 139] = tx_st_data          [ 273] ;
  assign tx_phy_preflop_1 [ 140] = tx_st_data          [ 274] ;
  assign tx_phy_preflop_1 [ 141] = tx_st_data          [ 275] ;
  assign tx_phy_preflop_1 [ 142] = tx_st_data          [ 276] ;
  assign tx_phy_preflop_1 [ 143] = tx_st_data          [ 277] ;
  assign tx_phy_preflop_1 [ 144] = tx_st_data          [ 278] ;
  assign tx_phy_preflop_1 [ 145] = tx_st_data          [ 279] ;
  assign tx_phy_preflop_1 [ 146] = tx_st_data          [ 280] ;
  assign tx_phy_preflop_1 [ 147] = tx_st_data          [ 281] ;
  assign tx_phy_preflop_1 [ 148] = tx_st_data          [ 282] ;
  assign tx_phy_preflop_1 [ 149] = tx_st_data          [ 283] ;
  assign tx_phy_preflop_1 [ 150] = tx_st_data          [ 284] ;
  assign tx_phy_preflop_1 [ 151] = tx_st_data          [ 285] ;
  assign tx_phy_preflop_1 [ 152] = tx_st_data          [ 286] ;
  assign tx_phy_preflop_1 [ 153] = tx_st_data          [ 287] ;
  assign tx_phy_preflop_1 [ 154] = tx_st_data          [ 288] ;
  assign tx_phy_preflop_1 [ 155] = tx_st_data          [ 289] ;
  assign tx_phy_preflop_1 [ 156] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 157] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 158] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 159] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 160] = tx_mrk_userbit[2]          ; // MARKER
  assign tx_phy_preflop_0 [ 161] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_0 [ 162] = tx_st_pushbit_r2           ;
  assign tx_phy_preflop_0 [ 163] = tx_st_data          [ 290] ;
  assign tx_phy_preflop_0 [ 164] = tx_st_data          [ 291] ;
  assign tx_phy_preflop_0 [ 165] = tx_st_data          [ 292] ;
  assign tx_phy_preflop_0 [ 166] = tx_st_data          [ 293] ;
  assign tx_phy_preflop_0 [ 167] = tx_st_data          [ 294] ;
  assign tx_phy_preflop_0 [ 168] = tx_st_data          [ 295] ;
  assign tx_phy_preflop_0 [ 169] = tx_st_data          [ 296] ;
  assign tx_phy_preflop_0 [ 170] = tx_st_data          [ 297] ;
  assign tx_phy_preflop_0 [ 171] = tx_st_data          [ 298] ;
  assign tx_phy_preflop_0 [ 172] = tx_st_data          [ 299] ;
  assign tx_phy_preflop_0 [ 173] = tx_st_data          [ 300] ;
  assign tx_phy_preflop_0 [ 174] = tx_st_data          [ 301] ;
  assign tx_phy_preflop_0 [ 175] = tx_st_data          [ 302] ;
  assign tx_phy_preflop_0 [ 176] = tx_st_data          [ 303] ;
  assign tx_phy_preflop_0 [ 177] = tx_st_data          [ 304] ;
  assign tx_phy_preflop_0 [ 178] = tx_st_data          [ 305] ;
  assign tx_phy_preflop_0 [ 179] = tx_st_data          [ 306] ;
  assign tx_phy_preflop_0 [ 180] = tx_st_data          [ 307] ;
  assign tx_phy_preflop_0 [ 181] = tx_st_data          [ 308] ;
  assign tx_phy_preflop_0 [ 182] = tx_st_data          [ 309] ;
  assign tx_phy_preflop_0 [ 183] = tx_st_data          [ 310] ;
  assign tx_phy_preflop_0 [ 184] = tx_st_data          [ 311] ;
  assign tx_phy_preflop_0 [ 185] = tx_st_data          [ 312] ;
  assign tx_phy_preflop_0 [ 186] = tx_st_data          [ 313] ;
  assign tx_phy_preflop_0 [ 187] = tx_st_data          [ 314] ;
  assign tx_phy_preflop_0 [ 188] = tx_st_data          [ 315] ;
  assign tx_phy_preflop_0 [ 189] = tx_st_data          [ 316] ;
  assign tx_phy_preflop_0 [ 190] = tx_st_data          [ 317] ;
  assign tx_phy_preflop_0 [ 191] = tx_st_data          [ 318] ;
  assign tx_phy_preflop_0 [ 192] = tx_st_data          [ 319] ;
  assign tx_phy_preflop_0 [ 193] = tx_st_data          [ 320] ;
  assign tx_phy_preflop_0 [ 194] = tx_st_data          [ 321] ;
  assign tx_phy_preflop_0 [ 195] = tx_st_data          [ 322] ;
  assign tx_phy_preflop_0 [ 196] = tx_st_data          [ 323] ;
  assign tx_phy_preflop_0 [ 197] = tx_st_data          [ 324] ;
  assign tx_phy_preflop_0 [ 198] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 199] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 200] = tx_st_data          [ 325] ;
  assign tx_phy_preflop_0 [ 201] = tx_st_data          [ 326] ;
  assign tx_phy_preflop_0 [ 202] = tx_st_data          [ 327] ;
  assign tx_phy_preflop_0 [ 203] = tx_st_data          [ 328] ;
  assign tx_phy_preflop_0 [ 204] = tx_st_data          [ 329] ;
  assign tx_phy_preflop_0 [ 205] = tx_st_data          [ 330] ;
  assign tx_phy_preflop_0 [ 206] = tx_st_data          [ 331] ;
  assign tx_phy_preflop_0 [ 207] = tx_st_data          [ 332] ;
  assign tx_phy_preflop_0 [ 208] = tx_st_data          [ 333] ;
  assign tx_phy_preflop_0 [ 209] = tx_st_data          [ 334] ;
  assign tx_phy_preflop_0 [ 210] = tx_st_data          [ 335] ;
  assign tx_phy_preflop_0 [ 211] = tx_st_data          [ 336] ;
  assign tx_phy_preflop_0 [ 212] = tx_st_data          [ 337] ;
  assign tx_phy_preflop_0 [ 213] = tx_st_data          [ 338] ;
  assign tx_phy_preflop_0 [ 214] = tx_st_data          [ 339] ;
  assign tx_phy_preflop_0 [ 215] = tx_st_data          [ 340] ;
  assign tx_phy_preflop_0 [ 216] = tx_st_data          [ 341] ;
  assign tx_phy_preflop_0 [ 217] = tx_st_data          [ 342] ;
  assign tx_phy_preflop_0 [ 218] = tx_st_data          [ 343] ;
  assign tx_phy_preflop_0 [ 219] = tx_st_data          [ 344] ;
  assign tx_phy_preflop_0 [ 220] = tx_st_data          [ 345] ;
  assign tx_phy_preflop_0 [ 221] = tx_st_data          [ 346] ;
  assign tx_phy_preflop_0 [ 222] = tx_st_data          [ 347] ;
  assign tx_phy_preflop_0 [ 223] = tx_st_data          [ 348] ;
  assign tx_phy_preflop_0 [ 224] = tx_st_data          [ 349] ;
  assign tx_phy_preflop_0 [ 225] = tx_st_data          [ 350] ;
  assign tx_phy_preflop_0 [ 226] = tx_st_data          [ 351] ;
  assign tx_phy_preflop_0 [ 227] = tx_st_data          [ 352] ;
  assign tx_phy_preflop_0 [ 228] = tx_st_data          [ 353] ;
  assign tx_phy_preflop_0 [ 229] = tx_st_data          [ 354] ;
  assign tx_phy_preflop_0 [ 230] = tx_st_data          [ 355] ;
  assign tx_phy_preflop_0 [ 231] = tx_st_data          [ 356] ;
  assign tx_phy_preflop_0 [ 232] = tx_st_data          [ 357] ;
  assign tx_phy_preflop_0 [ 233] = tx_st_data          [ 358] ;
  assign tx_phy_preflop_0 [ 234] = tx_st_data          [ 359] ;
  assign tx_phy_preflop_0 [ 235] = tx_st_data          [ 360] ;
  assign tx_phy_preflop_0 [ 236] = tx_st_data          [ 361] ;
  assign tx_phy_preflop_0 [ 237] = tx_st_data          [ 362] ;
  assign tx_phy_preflop_0 [ 238] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 239] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 160] = tx_mrk_userbit[2]          ; // MARKER
  assign tx_phy_preflop_1 [ 161] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_1 [ 162] = tx_st_data          [ 363] ;
  assign tx_phy_preflop_1 [ 163] = tx_st_data          [ 364] ;
  assign tx_phy_preflop_1 [ 164] = tx_st_data          [ 365] ;
  assign tx_phy_preflop_1 [ 165] = tx_st_data          [ 366] ;
  assign tx_phy_preflop_1 [ 166] = tx_st_data          [ 367] ;
  assign tx_phy_preflop_1 [ 167] = tx_st_data          [ 368] ;
  assign tx_phy_preflop_1 [ 168] = tx_st_data          [ 369] ;
  assign tx_phy_preflop_1 [ 169] = tx_st_data          [ 370] ;
  assign tx_phy_preflop_1 [ 170] = tx_st_data          [ 371] ;
  assign tx_phy_preflop_1 [ 171] = tx_st_data          [ 372] ;
  assign tx_phy_preflop_1 [ 172] = tx_st_data          [ 373] ;
  assign tx_phy_preflop_1 [ 173] = tx_st_data          [ 374] ;
  assign tx_phy_preflop_1 [ 174] = tx_st_data          [ 375] ;
  assign tx_phy_preflop_1 [ 175] = tx_st_data          [ 376] ;
  assign tx_phy_preflop_1 [ 176] = tx_st_data          [ 377] ;
  assign tx_phy_preflop_1 [ 177] = tx_st_data          [ 378] ;
  assign tx_phy_preflop_1 [ 178] = tx_st_data          [ 379] ;
  assign tx_phy_preflop_1 [ 179] = tx_st_data          [ 380] ;
  assign tx_phy_preflop_1 [ 180] = tx_st_data          [ 381] ;
  assign tx_phy_preflop_1 [ 181] = tx_st_data          [ 382] ;
  assign tx_phy_preflop_1 [ 182] = tx_st_data          [ 383] ;
  assign tx_phy_preflop_1 [ 183] = tx_st_data          [ 384] ;
  assign tx_phy_preflop_1 [ 184] = tx_st_data          [ 385] ;
  assign tx_phy_preflop_1 [ 185] = tx_st_data          [ 386] ;
  assign tx_phy_preflop_1 [ 186] = tx_st_data          [ 387] ;
  assign tx_phy_preflop_1 [ 187] = tx_st_data          [ 388] ;
  assign tx_phy_preflop_1 [ 188] = tx_st_data          [ 389] ;
  assign tx_phy_preflop_1 [ 189] = tx_st_data          [ 390] ;
  assign tx_phy_preflop_1 [ 190] = tx_st_data          [ 391] ;
  assign tx_phy_preflop_1 [ 191] = tx_st_data          [ 392] ;
  assign tx_phy_preflop_1 [ 192] = tx_st_data          [ 393] ;
  assign tx_phy_preflop_1 [ 193] = tx_st_data          [ 394] ;
  assign tx_phy_preflop_1 [ 194] = tx_st_data          [ 395] ;
  assign tx_phy_preflop_1 [ 195] = tx_st_data          [ 396] ;
  assign tx_phy_preflop_1 [ 196] = tx_st_data          [ 397] ;
  assign tx_phy_preflop_1 [ 197] = tx_st_data          [ 398] ;
  assign tx_phy_preflop_1 [ 198] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 199] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 200] = tx_st_data          [ 399] ;
  assign tx_phy_preflop_1 [ 201] = tx_st_data          [ 400] ;
  assign tx_phy_preflop_1 [ 202] = tx_st_data          [ 401] ;
  assign tx_phy_preflop_1 [ 203] = tx_st_data          [ 402] ;
  assign tx_phy_preflop_1 [ 204] = tx_st_data          [ 403] ;
  assign tx_phy_preflop_1 [ 205] = tx_st_data          [ 404] ;
  assign tx_phy_preflop_1 [ 206] = tx_st_data          [ 405] ;
  assign tx_phy_preflop_1 [ 207] = tx_st_data          [ 406] ;
  assign tx_phy_preflop_1 [ 208] = tx_st_data          [ 407] ;
  assign tx_phy_preflop_1 [ 209] = tx_st_data          [ 408] ;
  assign tx_phy_preflop_1 [ 210] = tx_st_data          [ 409] ;
  assign tx_phy_preflop_1 [ 211] = tx_st_data          [ 410] ;
  assign tx_phy_preflop_1 [ 212] = tx_st_data          [ 411] ;
  assign tx_phy_preflop_1 [ 213] = tx_st_data          [ 412] ;
  assign tx_phy_preflop_1 [ 214] = tx_st_data          [ 413] ;
  assign tx_phy_preflop_1 [ 215] = tx_st_data          [ 414] ;
  assign tx_phy_preflop_1 [ 216] = tx_st_data          [ 415] ;
  assign tx_phy_preflop_1 [ 217] = tx_st_data          [ 416] ;
  assign tx_phy_preflop_1 [ 218] = tx_st_data          [ 417] ;
  assign tx_phy_preflop_1 [ 219] = tx_st_data          [ 418] ;
  assign tx_phy_preflop_1 [ 220] = tx_st_data          [ 419] ;
  assign tx_phy_preflop_1 [ 221] = tx_st_data          [ 420] ;
  assign tx_phy_preflop_1 [ 222] = tx_st_data          [ 421] ;
  assign tx_phy_preflop_1 [ 223] = tx_st_data          [ 422] ;
  assign tx_phy_preflop_1 [ 224] = tx_st_data          [ 423] ;
  assign tx_phy_preflop_1 [ 225] = tx_st_data          [ 424] ;
  assign tx_phy_preflop_1 [ 226] = tx_st_data          [ 425] ;
  assign tx_phy_preflop_1 [ 227] = tx_st_data          [ 426] ;
  assign tx_phy_preflop_1 [ 228] = tx_st_data          [ 427] ;
  assign tx_phy_preflop_1 [ 229] = tx_st_data          [ 428] ;
  assign tx_phy_preflop_1 [ 230] = tx_st_data          [ 429] ;
  assign tx_phy_preflop_1 [ 231] = tx_st_data          [ 430] ;
  assign tx_phy_preflop_1 [ 232] = tx_st_data          [ 431] ;
  assign tx_phy_preflop_1 [ 233] = tx_st_data          [ 432] ;
  assign tx_phy_preflop_1 [ 234] = tx_st_data          [ 433] ;
  assign tx_phy_preflop_1 [ 235] = tx_st_data          [ 434] ;
  assign tx_phy_preflop_1 [ 236] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 237] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 238] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 239] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 240] = tx_mrk_userbit[3]          ; // MARKER
  assign tx_phy_preflop_0 [ 241] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_0 [ 242] = tx_st_pushbit_r3           ;
  assign tx_phy_preflop_0 [ 243] = tx_st_data          [ 435] ;
  assign tx_phy_preflop_0 [ 244] = tx_st_data          [ 436] ;
  assign tx_phy_preflop_0 [ 245] = tx_st_data          [ 437] ;
  assign tx_phy_preflop_0 [ 246] = tx_st_data          [ 438] ;
  assign tx_phy_preflop_0 [ 247] = tx_st_data          [ 439] ;
  assign tx_phy_preflop_0 [ 248] = tx_st_data          [ 440] ;
  assign tx_phy_preflop_0 [ 249] = tx_st_data          [ 441] ;
  assign tx_phy_preflop_0 [ 250] = tx_st_data          [ 442] ;
  assign tx_phy_preflop_0 [ 251] = tx_st_data          [ 443] ;
  assign tx_phy_preflop_0 [ 252] = tx_st_data          [ 444] ;
  assign tx_phy_preflop_0 [ 253] = tx_st_data          [ 445] ;
  assign tx_phy_preflop_0 [ 254] = tx_st_data          [ 446] ;
  assign tx_phy_preflop_0 [ 255] = tx_st_data          [ 447] ;
  assign tx_phy_preflop_0 [ 256] = tx_st_data          [ 448] ;
  assign tx_phy_preflop_0 [ 257] = tx_st_data          [ 449] ;
  assign tx_phy_preflop_0 [ 258] = tx_st_data          [ 450] ;
  assign tx_phy_preflop_0 [ 259] = tx_st_data          [ 451] ;
  assign tx_phy_preflop_0 [ 260] = tx_st_data          [ 452] ;
  assign tx_phy_preflop_0 [ 261] = tx_st_data          [ 453] ;
  assign tx_phy_preflop_0 [ 262] = tx_st_data          [ 454] ;
  assign tx_phy_preflop_0 [ 263] = tx_st_data          [ 455] ;
  assign tx_phy_preflop_0 [ 264] = tx_st_data          [ 456] ;
  assign tx_phy_preflop_0 [ 265] = tx_st_data          [ 457] ;
  assign tx_phy_preflop_0 [ 266] = tx_st_data          [ 458] ;
  assign tx_phy_preflop_0 [ 267] = tx_st_data          [ 459] ;
  assign tx_phy_preflop_0 [ 268] = tx_st_data          [ 460] ;
  assign tx_phy_preflop_0 [ 269] = tx_st_data          [ 461] ;
  assign tx_phy_preflop_0 [ 270] = tx_st_data          [ 462] ;
  assign tx_phy_preflop_0 [ 271] = tx_st_data          [ 463] ;
  assign tx_phy_preflop_0 [ 272] = tx_st_data          [ 464] ;
  assign tx_phy_preflop_0 [ 273] = tx_st_data          [ 465] ;
  assign tx_phy_preflop_0 [ 274] = tx_st_data          [ 466] ;
  assign tx_phy_preflop_0 [ 275] = tx_st_data          [ 467] ;
  assign tx_phy_preflop_0 [ 276] = tx_st_data          [ 468] ;
  assign tx_phy_preflop_0 [ 277] = tx_st_data          [ 469] ;
  assign tx_phy_preflop_0 [ 278] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 279] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 280] = tx_st_data          [ 470] ;
  assign tx_phy_preflop_0 [ 281] = tx_st_data          [ 471] ;
  assign tx_phy_preflop_0 [ 282] = tx_st_data          [ 472] ;
  assign tx_phy_preflop_0 [ 283] = tx_st_data          [ 473] ;
  assign tx_phy_preflop_0 [ 284] = tx_st_data          [ 474] ;
  assign tx_phy_preflop_0 [ 285] = tx_st_data          [ 475] ;
  assign tx_phy_preflop_0 [ 286] = tx_st_data          [ 476] ;
  assign tx_phy_preflop_0 [ 287] = tx_st_data          [ 477] ;
  assign tx_phy_preflop_0 [ 288] = tx_st_data          [ 478] ;
  assign tx_phy_preflop_0 [ 289] = tx_st_data          [ 479] ;
  assign tx_phy_preflop_0 [ 290] = tx_st_data          [ 480] ;
  assign tx_phy_preflop_0 [ 291] = tx_st_data          [ 481] ;
  assign tx_phy_preflop_0 [ 292] = tx_st_data          [ 482] ;
  assign tx_phy_preflop_0 [ 293] = tx_st_data          [ 483] ;
  assign tx_phy_preflop_0 [ 294] = tx_st_data          [ 484] ;
  assign tx_phy_preflop_0 [ 295] = tx_st_data          [ 485] ;
  assign tx_phy_preflop_0 [ 296] = tx_st_data          [ 486] ;
  assign tx_phy_preflop_0 [ 297] = tx_st_data          [ 487] ;
  assign tx_phy_preflop_0 [ 298] = tx_st_data          [ 488] ;
  assign tx_phy_preflop_0 [ 299] = tx_st_data          [ 489] ;
  assign tx_phy_preflop_0 [ 300] = tx_st_data          [ 490] ;
  assign tx_phy_preflop_0 [ 301] = tx_st_data          [ 491] ;
  assign tx_phy_preflop_0 [ 302] = tx_st_data          [ 492] ;
  assign tx_phy_preflop_0 [ 303] = tx_st_data          [ 493] ;
  assign tx_phy_preflop_0 [ 304] = tx_st_data          [ 494] ;
  assign tx_phy_preflop_0 [ 305] = tx_st_data          [ 495] ;
  assign tx_phy_preflop_0 [ 306] = tx_st_data          [ 496] ;
  assign tx_phy_preflop_0 [ 307] = tx_st_data          [ 497] ;
  assign tx_phy_preflop_0 [ 308] = tx_st_data          [ 498] ;
  assign tx_phy_preflop_0 [ 309] = tx_st_data          [ 499] ;
  assign tx_phy_preflop_0 [ 310] = tx_st_data          [ 500] ;
  assign tx_phy_preflop_0 [ 311] = tx_st_data          [ 501] ;
  assign tx_phy_preflop_0 [ 312] = tx_st_data          [ 502] ;
  assign tx_phy_preflop_0 [ 313] = tx_st_data          [ 503] ;
  assign tx_phy_preflop_0 [ 314] = tx_st_data          [ 504] ;
  assign tx_phy_preflop_0 [ 315] = tx_st_data          [ 505] ;
  assign tx_phy_preflop_0 [ 316] = tx_st_data          [ 506] ;
  assign tx_phy_preflop_0 [ 317] = tx_st_data          [ 507] ;
  assign tx_phy_preflop_0 [ 318] = 1'b0                       ; // DBI
  assign tx_phy_preflop_0 [ 319] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 240] = tx_mrk_userbit[3]          ; // MARKER
  assign tx_phy_preflop_1 [ 241] = 1'b0                       ; // STROBE (unused)
  assign tx_phy_preflop_1 [ 242] = tx_st_data          [ 508] ;
  assign tx_phy_preflop_1 [ 243] = tx_st_data          [ 509] ;
  assign tx_phy_preflop_1 [ 244] = tx_st_data          [ 510] ;
  assign tx_phy_preflop_1 [ 245] = tx_st_data          [ 511] ;
  assign tx_phy_preflop_1 [ 246] = tx_st_data          [ 512] ;
  assign tx_phy_preflop_1 [ 247] = tx_st_data          [ 513] ;
  assign tx_phy_preflop_1 [ 248] = tx_st_data          [ 514] ;
  assign tx_phy_preflop_1 [ 249] = tx_st_data          [ 515] ;
  assign tx_phy_preflop_1 [ 250] = tx_st_data          [ 516] ;
  assign tx_phy_preflop_1 [ 251] = tx_st_data          [ 517] ;
  assign tx_phy_preflop_1 [ 252] = tx_st_data          [ 518] ;
  assign tx_phy_preflop_1 [ 253] = tx_st_data          [ 519] ;
  assign tx_phy_preflop_1 [ 254] = tx_st_data          [ 520] ;
  assign tx_phy_preflop_1 [ 255] = tx_st_data          [ 521] ;
  assign tx_phy_preflop_1 [ 256] = tx_st_data          [ 522] ;
  assign tx_phy_preflop_1 [ 257] = tx_st_data          [ 523] ;
  assign tx_phy_preflop_1 [ 258] = tx_st_data          [ 524] ;
  assign tx_phy_preflop_1 [ 259] = tx_st_data          [ 525] ;
  assign tx_phy_preflop_1 [ 260] = tx_st_data          [ 526] ;
  assign tx_phy_preflop_1 [ 261] = tx_st_data          [ 527] ;
  assign tx_phy_preflop_1 [ 262] = tx_st_data          [ 528] ;
  assign tx_phy_preflop_1 [ 263] = tx_st_data          [ 529] ;
  assign tx_phy_preflop_1 [ 264] = tx_st_data          [ 530] ;
  assign tx_phy_preflop_1 [ 265] = tx_st_data          [ 531] ;
  assign tx_phy_preflop_1 [ 266] = tx_st_data          [ 532] ;
  assign tx_phy_preflop_1 [ 267] = tx_st_data          [ 533] ;
  assign tx_phy_preflop_1 [ 268] = tx_st_data          [ 534] ;
  assign tx_phy_preflop_1 [ 269] = tx_st_data          [ 535] ;
  assign tx_phy_preflop_1 [ 270] = tx_st_data          [ 536] ;
  assign tx_phy_preflop_1 [ 271] = tx_st_data          [ 537] ;
  assign tx_phy_preflop_1 [ 272] = tx_st_data          [ 538] ;
  assign tx_phy_preflop_1 [ 273] = tx_st_data          [ 539] ;
  assign tx_phy_preflop_1 [ 274] = tx_st_data          [ 540] ;
  assign tx_phy_preflop_1 [ 275] = tx_st_data          [ 541] ;
  assign tx_phy_preflop_1 [ 276] = tx_st_data          [ 542] ;
  assign tx_phy_preflop_1 [ 277] = tx_st_data          [ 543] ;
  assign tx_phy_preflop_1 [ 278] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 279] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 280] = tx_st_data          [ 544] ;
  assign tx_phy_preflop_1 [ 281] = tx_st_data          [ 545] ;
  assign tx_phy_preflop_1 [ 282] = tx_st_data          [ 546] ;
  assign tx_phy_preflop_1 [ 283] = tx_st_data          [ 547] ;
  assign tx_phy_preflop_1 [ 284] = tx_st_data          [ 548] ;
  assign tx_phy_preflop_1 [ 285] = tx_st_data          [ 549] ;
  assign tx_phy_preflop_1 [ 286] = tx_st_data          [ 550] ;
  assign tx_phy_preflop_1 [ 287] = tx_st_data          [ 551] ;
  assign tx_phy_preflop_1 [ 288] = tx_st_data          [ 552] ;
  assign tx_phy_preflop_1 [ 289] = tx_st_data          [ 553] ;
  assign tx_phy_preflop_1 [ 290] = tx_st_data          [ 554] ;
  assign tx_phy_preflop_1 [ 291] = tx_st_data          [ 555] ;
  assign tx_phy_preflop_1 [ 292] = tx_st_data          [ 556] ;
  assign tx_phy_preflop_1 [ 293] = tx_st_data          [ 557] ;
  assign tx_phy_preflop_1 [ 294] = tx_st_data          [ 558] ;
  assign tx_phy_preflop_1 [ 295] = tx_st_data          [ 559] ;
  assign tx_phy_preflop_1 [ 296] = tx_st_data          [ 560] ;
  assign tx_phy_preflop_1 [ 297] = tx_st_data          [ 561] ;
  assign tx_phy_preflop_1 [ 298] = tx_st_data          [ 562] ;
  assign tx_phy_preflop_1 [ 299] = tx_st_data          [ 563] ;
  assign tx_phy_preflop_1 [ 300] = tx_st_data          [ 564] ;
  assign tx_phy_preflop_1 [ 301] = tx_st_data          [ 565] ;
  assign tx_phy_preflop_1 [ 302] = tx_st_data          [ 566] ;
  assign tx_phy_preflop_1 [ 303] = tx_st_data          [ 567] ;
  assign tx_phy_preflop_1 [ 304] = tx_st_data          [ 568] ;
  assign tx_phy_preflop_1 [ 305] = tx_st_data          [ 569] ;
  assign tx_phy_preflop_1 [ 306] = tx_st_data          [ 570] ;
  assign tx_phy_preflop_1 [ 307] = tx_st_data          [ 571] ;
  assign tx_phy_preflop_1 [ 308] = tx_st_data          [ 572] ;
  assign tx_phy_preflop_1 [ 309] = tx_st_data          [ 573] ;
  assign tx_phy_preflop_1 [ 310] = tx_st_data          [ 574] ;
  assign tx_phy_preflop_1 [ 311] = tx_st_data          [ 575] ;
  assign tx_phy_preflop_1 [ 312] = tx_st_data          [ 576] ;
  assign tx_phy_preflop_1 [ 313] = tx_st_data          [ 577] ;
  assign tx_phy_preflop_1 [ 314] = tx_st_data          [ 578] ;
  assign tx_phy_preflop_1 [ 315] = tx_st_data          [ 579] ;
  assign tx_phy_preflop_1 [ 316] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 317] = 1'b0                       ;
  assign tx_phy_preflop_1 [ 318] = 1'b0                       ; // DBI
  assign tx_phy_preflop_1 [ 319] = 1'b0                       ; // DBI
// TX Section
//////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////
// RX Section

//   RX_CH_WIDTH           = 320; // Gen2Only running at Quarter Rate
//   RX_DATA_WIDTH         = 296; // Usable Data per Channel
//   RX_PERSISTENT_STROBE  = 1'b1;
//   RX_PERSISTENT_MARKER  = 1'b1;
//   RX_STROBE_GEN2_LOC    = 'd1;
//   RX_MARKER_GEN2_LOC    = 'd0;
//   RX_STROBE_GEN1_LOC    = 'd38;
//   RX_MARKER_GEN1_LOC    = 'd39;
//   RX_ENABLE_STROBE      = 1'b1;
//   RX_ENABLE_MARKER      = 1'b1;
//   RX_DBI_PRESENT        = 1'b1;
//   RX_REG_PHY            = 1'b0;

  localparam RX_REG_PHY    = 1'b0;  // If set, this enables boundary FF for timing reasons

  logic [ 319:   0]                              rx_phy_postflop_0             ;
  logic [ 319:   0]                              rx_phy_postflop_1             ;
  logic [ 319:   0]                              rx_phy_flop_0_reg             ;
  logic [ 319:   0]                              rx_phy_flop_1_reg             ;

  always_ff @(posedge clk_rd or negedge rst_rd_n)
  if (~rst_rd_n)
  begin
    rx_phy_flop_0_reg                       <= 320'b0                                  ;
    rx_phy_flop_1_reg                       <= 320'b0                                  ;
  end
  else
  begin
    rx_phy_flop_0_reg                       <= rx_phy0                                 ;
    rx_phy_flop_1_reg                       <= rx_phy1                                 ;
  end


  assign rx_phy_postflop_0                  = RX_REG_PHY ? rx_phy_flop_0_reg : rx_phy0               ;
  assign rx_phy_postflop_1                  = RX_REG_PHY ? rx_phy_flop_1_reg : rx_phy1               ;

  logic                                          rx_st_credit_r0               ;
  logic                                          rx_st_credit_r1               ;
  logic                                          rx_st_credit_r2               ;
  logic                                          rx_st_credit_r3               ;

  // Asymmetric Credit Logic
  assign rx_st_credit         [   0 +:   1] = rx_st_credit_r0                    ;
  assign rx_st_credit         [   1 +:   1] = rx_st_credit_r1                    ;
  assign rx_st_credit         [   2 +:   1] = rx_st_credit_r2                    ;
  assign rx_st_credit         [   3 +:   1] = rx_st_credit_r3                    ;

//       MARKER                     = rx_phy_postflop_0 [   0]
//       STROBE                     = rx_phy_postflop_0 [   1]
  assign rx_st_credit_r0            = rx_phy_postflop_0 [   2];
//       nc                         = rx_phy_postflop_0 [   3];
//       nc                         = rx_phy_postflop_0 [   4];
//       nc                         = rx_phy_postflop_0 [   5];
//       nc                         = rx_phy_postflop_0 [   6];
//       nc                         = rx_phy_postflop_0 [   7];
//       nc                         = rx_phy_postflop_0 [   8];
//       nc                         = rx_phy_postflop_0 [   9];
//       nc                         = rx_phy_postflop_0 [  10];
//       nc                         = rx_phy_postflop_0 [  11];
//       nc                         = rx_phy_postflop_0 [  12];
//       nc                         = rx_phy_postflop_0 [  13];
//       nc                         = rx_phy_postflop_0 [  14];
//       nc                         = rx_phy_postflop_0 [  15];
//       nc                         = rx_phy_postflop_0 [  16];
//       nc                         = rx_phy_postflop_0 [  17];
//       nc                         = rx_phy_postflop_0 [  18];
//       nc                         = rx_phy_postflop_0 [  19];
//       nc                         = rx_phy_postflop_0 [  20];
//       nc                         = rx_phy_postflop_0 [  21];
//       nc                         = rx_phy_postflop_0 [  22];
//       nc                         = rx_phy_postflop_0 [  23];
//       nc                         = rx_phy_postflop_0 [  24];
//       nc                         = rx_phy_postflop_0 [  25];
//       nc                         = rx_phy_postflop_0 [  26];
//       nc                         = rx_phy_postflop_0 [  27];
//       nc                         = rx_phy_postflop_0 [  28];
//       nc                         = rx_phy_postflop_0 [  29];
//       nc                         = rx_phy_postflop_0 [  30];
//       nc                         = rx_phy_postflop_0 [  31];
//       nc                         = rx_phy_postflop_0 [  32];
//       nc                         = rx_phy_postflop_0 [  33];
//       nc                         = rx_phy_postflop_0 [  34];
//       nc                         = rx_phy_postflop_0 [  35];
//       nc                         = rx_phy_postflop_0 [  36];
//       nc                         = rx_phy_postflop_0 [  37];
//       DBI                        = rx_phy_postflop_0 [  38];
//       DBI                        = rx_phy_postflop_0 [  39];
//       nc                         = rx_phy_postflop_0 [  40];
//       nc                         = rx_phy_postflop_0 [  41];
//       nc                         = rx_phy_postflop_0 [  42];
//       nc                         = rx_phy_postflop_0 [  43];
//       nc                         = rx_phy_postflop_0 [  44];
//       nc                         = rx_phy_postflop_0 [  45];
//       nc                         = rx_phy_postflop_0 [  46];
//       nc                         = rx_phy_postflop_0 [  47];
//       nc                         = rx_phy_postflop_0 [  48];
//       nc                         = rx_phy_postflop_0 [  49];
//       nc                         = rx_phy_postflop_0 [  50];
//       nc                         = rx_phy_postflop_0 [  51];
//       nc                         = rx_phy_postflop_0 [  52];
//       nc                         = rx_phy_postflop_0 [  53];
//       nc                         = rx_phy_postflop_0 [  54];
//       nc                         = rx_phy_postflop_0 [  55];
//       nc                         = rx_phy_postflop_0 [  56];
//       nc                         = rx_phy_postflop_0 [  57];
//       nc                         = rx_phy_postflop_0 [  58];
//       nc                         = rx_phy_postflop_0 [  59];
//       nc                         = rx_phy_postflop_0 [  60];
//       nc                         = rx_phy_postflop_0 [  61];
//       nc                         = rx_phy_postflop_0 [  62];
//       nc                         = rx_phy_postflop_0 [  63];
//       nc                         = rx_phy_postflop_0 [  64];
//       nc                         = rx_phy_postflop_0 [  65];
//       nc                         = rx_phy_postflop_0 [  66];
//       nc                         = rx_phy_postflop_0 [  67];
//       nc                         = rx_phy_postflop_0 [  68];
//       nc                         = rx_phy_postflop_0 [  69];
//       nc                         = rx_phy_postflop_0 [  70];
//       nc                         = rx_phy_postflop_0 [  71];
//       nc                         = rx_phy_postflop_0 [  72];
//       nc                         = rx_phy_postflop_0 [  73];
//       nc                         = rx_phy_postflop_0 [  74];
//       nc                         = rx_phy_postflop_0 [  75];
//       nc                         = rx_phy_postflop_0 [  76];
//       nc                         = rx_phy_postflop_0 [  77];
//       DBI                        = rx_phy_postflop_0 [  78];
//       DBI                        = rx_phy_postflop_0 [  79];
//       MARKER                     = rx_phy_postflop_1 [   0]
//       STROBE                     = rx_phy_postflop_1 [   1]
//       nc                         = rx_phy_postflop_1 [   2];
//       nc                         = rx_phy_postflop_1 [   3];
//       nc                         = rx_phy_postflop_1 [   4];
//       nc                         = rx_phy_postflop_1 [   5];
//       nc                         = rx_phy_postflop_1 [   6];
//       nc                         = rx_phy_postflop_1 [   7];
//       nc                         = rx_phy_postflop_1 [   8];
//       nc                         = rx_phy_postflop_1 [   9];
//       nc                         = rx_phy_postflop_1 [  10];
//       nc                         = rx_phy_postflop_1 [  11];
//       nc                         = rx_phy_postflop_1 [  12];
//       nc                         = rx_phy_postflop_1 [  13];
//       nc                         = rx_phy_postflop_1 [  14];
//       nc                         = rx_phy_postflop_1 [  15];
//       nc                         = rx_phy_postflop_1 [  16];
//       nc                         = rx_phy_postflop_1 [  17];
//       nc                         = rx_phy_postflop_1 [  18];
//       nc                         = rx_phy_postflop_1 [  19];
//       nc                         = rx_phy_postflop_1 [  20];
//       nc                         = rx_phy_postflop_1 [  21];
//       nc                         = rx_phy_postflop_1 [  22];
//       nc                         = rx_phy_postflop_1 [  23];
//       nc                         = rx_phy_postflop_1 [  24];
//       nc                         = rx_phy_postflop_1 [  25];
//       nc                         = rx_phy_postflop_1 [  26];
//       nc                         = rx_phy_postflop_1 [  27];
//       nc                         = rx_phy_postflop_1 [  28];
//       nc                         = rx_phy_postflop_1 [  29];
//       nc                         = rx_phy_postflop_1 [  30];
//       nc                         = rx_phy_postflop_1 [  31];
//       nc                         = rx_phy_postflop_1 [  32];
//       nc                         = rx_phy_postflop_1 [  33];
//       nc                         = rx_phy_postflop_1 [  34];
//       nc                         = rx_phy_postflop_1 [  35];
//       nc                         = rx_phy_postflop_1 [  36];
//       nc                         = rx_phy_postflop_1 [  37];
//       DBI                        = rx_phy_postflop_1 [  38];
//       DBI                        = rx_phy_postflop_1 [  39];
//       nc                         = rx_phy_postflop_1 [  40];
//       nc                         = rx_phy_postflop_1 [  41];
//       nc                         = rx_phy_postflop_1 [  42];
//       nc                         = rx_phy_postflop_1 [  43];
//       nc                         = rx_phy_postflop_1 [  44];
//       nc                         = rx_phy_postflop_1 [  45];
//       nc                         = rx_phy_postflop_1 [  46];
//       nc                         = rx_phy_postflop_1 [  47];
//       nc                         = rx_phy_postflop_1 [  48];
//       nc                         = rx_phy_postflop_1 [  49];
//       nc                         = rx_phy_postflop_1 [  50];
//       nc                         = rx_phy_postflop_1 [  51];
//       nc                         = rx_phy_postflop_1 [  52];
//       nc                         = rx_phy_postflop_1 [  53];
//       nc                         = rx_phy_postflop_1 [  54];
//       nc                         = rx_phy_postflop_1 [  55];
//       nc                         = rx_phy_postflop_1 [  56];
//       nc                         = rx_phy_postflop_1 [  57];
//       nc                         = rx_phy_postflop_1 [  58];
//       nc                         = rx_phy_postflop_1 [  59];
//       nc                         = rx_phy_postflop_1 [  60];
//       nc                         = rx_phy_postflop_1 [  61];
//       nc                         = rx_phy_postflop_1 [  62];
//       nc                         = rx_phy_postflop_1 [  63];
//       nc                         = rx_phy_postflop_1 [  64];
//       nc                         = rx_phy_postflop_1 [  65];
//       nc                         = rx_phy_postflop_1 [  66];
//       nc                         = rx_phy_postflop_1 [  67];
//       nc                         = rx_phy_postflop_1 [  68];
//       nc                         = rx_phy_postflop_1 [  69];
//       nc                         = rx_phy_postflop_1 [  70];
//       nc                         = rx_phy_postflop_1 [  71];
//       nc                         = rx_phy_postflop_1 [  72];
//       nc                         = rx_phy_postflop_1 [  73];
//       nc                         = rx_phy_postflop_1 [  74];
//       nc                         = rx_phy_postflop_1 [  75];
//       nc                         = rx_phy_postflop_1 [  76];
//       nc                         = rx_phy_postflop_1 [  77];
//       DBI                        = rx_phy_postflop_1 [  78];
//       DBI                        = rx_phy_postflop_1 [  79];
//       MARKER                     = rx_phy_postflop_0 [  80]
//       STROBE                     = rx_phy_postflop_0 [  81]
  assign rx_st_credit_r1            = rx_phy_postflop_0 [  82];
//       nc                         = rx_phy_postflop_0 [  83];
//       nc                         = rx_phy_postflop_0 [  84];
//       nc                         = rx_phy_postflop_0 [  85];
//       nc                         = rx_phy_postflop_0 [  86];
//       nc                         = rx_phy_postflop_0 [  87];
//       nc                         = rx_phy_postflop_0 [  88];
//       nc                         = rx_phy_postflop_0 [  89];
//       nc                         = rx_phy_postflop_0 [  90];
//       nc                         = rx_phy_postflop_0 [  91];
//       nc                         = rx_phy_postflop_0 [  92];
//       nc                         = rx_phy_postflop_0 [  93];
//       nc                         = rx_phy_postflop_0 [  94];
//       nc                         = rx_phy_postflop_0 [  95];
//       nc                         = rx_phy_postflop_0 [  96];
//       nc                         = rx_phy_postflop_0 [  97];
//       nc                         = rx_phy_postflop_0 [  98];
//       nc                         = rx_phy_postflop_0 [  99];
//       nc                         = rx_phy_postflop_0 [ 100];
//       nc                         = rx_phy_postflop_0 [ 101];
//       nc                         = rx_phy_postflop_0 [ 102];
//       nc                         = rx_phy_postflop_0 [ 103];
//       nc                         = rx_phy_postflop_0 [ 104];
//       nc                         = rx_phy_postflop_0 [ 105];
//       nc                         = rx_phy_postflop_0 [ 106];
//       nc                         = rx_phy_postflop_0 [ 107];
//       nc                         = rx_phy_postflop_0 [ 108];
//       nc                         = rx_phy_postflop_0 [ 109];
//       nc                         = rx_phy_postflop_0 [ 110];
//       nc                         = rx_phy_postflop_0 [ 111];
//       nc                         = rx_phy_postflop_0 [ 112];
//       nc                         = rx_phy_postflop_0 [ 113];
//       nc                         = rx_phy_postflop_0 [ 114];
//       nc                         = rx_phy_postflop_0 [ 115];
//       nc                         = rx_phy_postflop_0 [ 116];
//       nc                         = rx_phy_postflop_0 [ 117];
//       DBI                        = rx_phy_postflop_0 [ 118];
//       DBI                        = rx_phy_postflop_0 [ 119];
//       nc                         = rx_phy_postflop_0 [ 120];
//       nc                         = rx_phy_postflop_0 [ 121];
//       nc                         = rx_phy_postflop_0 [ 122];
//       nc                         = rx_phy_postflop_0 [ 123];
//       nc                         = rx_phy_postflop_0 [ 124];
//       nc                         = rx_phy_postflop_0 [ 125];
//       nc                         = rx_phy_postflop_0 [ 126];
//       nc                         = rx_phy_postflop_0 [ 127];
//       nc                         = rx_phy_postflop_0 [ 128];
//       nc                         = rx_phy_postflop_0 [ 129];
//       nc                         = rx_phy_postflop_0 [ 130];
//       nc                         = rx_phy_postflop_0 [ 131];
//       nc                         = rx_phy_postflop_0 [ 132];
//       nc                         = rx_phy_postflop_0 [ 133];
//       nc                         = rx_phy_postflop_0 [ 134];
//       nc                         = rx_phy_postflop_0 [ 135];
//       nc                         = rx_phy_postflop_0 [ 136];
//       nc                         = rx_phy_postflop_0 [ 137];
//       nc                         = rx_phy_postflop_0 [ 138];
//       nc                         = rx_phy_postflop_0 [ 139];
//       nc                         = rx_phy_postflop_0 [ 140];
//       nc                         = rx_phy_postflop_0 [ 141];
//       nc                         = rx_phy_postflop_0 [ 142];
//       nc                         = rx_phy_postflop_0 [ 143];
//       nc                         = rx_phy_postflop_0 [ 144];
//       nc                         = rx_phy_postflop_0 [ 145];
//       nc                         = rx_phy_postflop_0 [ 146];
//       nc                         = rx_phy_postflop_0 [ 147];
//       nc                         = rx_phy_postflop_0 [ 148];
//       nc                         = rx_phy_postflop_0 [ 149];
//       nc                         = rx_phy_postflop_0 [ 150];
//       nc                         = rx_phy_postflop_0 [ 151];
//       nc                         = rx_phy_postflop_0 [ 152];
//       nc                         = rx_phy_postflop_0 [ 153];
//       nc                         = rx_phy_postflop_0 [ 154];
//       nc                         = rx_phy_postflop_0 [ 155];
//       nc                         = rx_phy_postflop_0 [ 156];
//       nc                         = rx_phy_postflop_0 [ 157];
//       DBI                        = rx_phy_postflop_0 [ 158];
//       DBI                        = rx_phy_postflop_0 [ 159];
//       MARKER                     = rx_phy_postflop_1 [  80]
//       STROBE                     = rx_phy_postflop_1 [  81]
//       nc                         = rx_phy_postflop_1 [  82];
//       nc                         = rx_phy_postflop_1 [  83];
//       nc                         = rx_phy_postflop_1 [  84];
//       nc                         = rx_phy_postflop_1 [  85];
//       nc                         = rx_phy_postflop_1 [  86];
//       nc                         = rx_phy_postflop_1 [  87];
//       nc                         = rx_phy_postflop_1 [  88];
//       nc                         = rx_phy_postflop_1 [  89];
//       nc                         = rx_phy_postflop_1 [  90];
//       nc                         = rx_phy_postflop_1 [  91];
//       nc                         = rx_phy_postflop_1 [  92];
//       nc                         = rx_phy_postflop_1 [  93];
//       nc                         = rx_phy_postflop_1 [  94];
//       nc                         = rx_phy_postflop_1 [  95];
//       nc                         = rx_phy_postflop_1 [  96];
//       nc                         = rx_phy_postflop_1 [  97];
//       nc                         = rx_phy_postflop_1 [  98];
//       nc                         = rx_phy_postflop_1 [  99];
//       nc                         = rx_phy_postflop_1 [ 100];
//       nc                         = rx_phy_postflop_1 [ 101];
//       nc                         = rx_phy_postflop_1 [ 102];
//       nc                         = rx_phy_postflop_1 [ 103];
//       nc                         = rx_phy_postflop_1 [ 104];
//       nc                         = rx_phy_postflop_1 [ 105];
//       nc                         = rx_phy_postflop_1 [ 106];
//       nc                         = rx_phy_postflop_1 [ 107];
//       nc                         = rx_phy_postflop_1 [ 108];
//       nc                         = rx_phy_postflop_1 [ 109];
//       nc                         = rx_phy_postflop_1 [ 110];
//       nc                         = rx_phy_postflop_1 [ 111];
//       nc                         = rx_phy_postflop_1 [ 112];
//       nc                         = rx_phy_postflop_1 [ 113];
//       nc                         = rx_phy_postflop_1 [ 114];
//       nc                         = rx_phy_postflop_1 [ 115];
//       nc                         = rx_phy_postflop_1 [ 116];
//       nc                         = rx_phy_postflop_1 [ 117];
//       DBI                        = rx_phy_postflop_1 [ 118];
//       DBI                        = rx_phy_postflop_1 [ 119];
//       nc                         = rx_phy_postflop_1 [ 120];
//       nc                         = rx_phy_postflop_1 [ 121];
//       nc                         = rx_phy_postflop_1 [ 122];
//       nc                         = rx_phy_postflop_1 [ 123];
//       nc                         = rx_phy_postflop_1 [ 124];
//       nc                         = rx_phy_postflop_1 [ 125];
//       nc                         = rx_phy_postflop_1 [ 126];
//       nc                         = rx_phy_postflop_1 [ 127];
//       nc                         = rx_phy_postflop_1 [ 128];
//       nc                         = rx_phy_postflop_1 [ 129];
//       nc                         = rx_phy_postflop_1 [ 130];
//       nc                         = rx_phy_postflop_1 [ 131];
//       nc                         = rx_phy_postflop_1 [ 132];
//       nc                         = rx_phy_postflop_1 [ 133];
//       nc                         = rx_phy_postflop_1 [ 134];
//       nc                         = rx_phy_postflop_1 [ 135];
//       nc                         = rx_phy_postflop_1 [ 136];
//       nc                         = rx_phy_postflop_1 [ 137];
//       nc                         = rx_phy_postflop_1 [ 138];
//       nc                         = rx_phy_postflop_1 [ 139];
//       nc                         = rx_phy_postflop_1 [ 140];
//       nc                         = rx_phy_postflop_1 [ 141];
//       nc                         = rx_phy_postflop_1 [ 142];
//       nc                         = rx_phy_postflop_1 [ 143];
//       nc                         = rx_phy_postflop_1 [ 144];
//       nc                         = rx_phy_postflop_1 [ 145];
//       nc                         = rx_phy_postflop_1 [ 146];
//       nc                         = rx_phy_postflop_1 [ 147];
//       nc                         = rx_phy_postflop_1 [ 148];
//       nc                         = rx_phy_postflop_1 [ 149];
//       nc                         = rx_phy_postflop_1 [ 150];
//       nc                         = rx_phy_postflop_1 [ 151];
//       nc                         = rx_phy_postflop_1 [ 152];
//       nc                         = rx_phy_postflop_1 [ 153];
//       nc                         = rx_phy_postflop_1 [ 154];
//       nc                         = rx_phy_postflop_1 [ 155];
//       nc                         = rx_phy_postflop_1 [ 156];
//       nc                         = rx_phy_postflop_1 [ 157];
//       DBI                        = rx_phy_postflop_1 [ 158];
//       DBI                        = rx_phy_postflop_1 [ 159];
//       MARKER                     = rx_phy_postflop_0 [ 160]
//       STROBE                     = rx_phy_postflop_0 [ 161]
  assign rx_st_credit_r2            = rx_phy_postflop_0 [ 162];
//       nc                         = rx_phy_postflop_0 [ 163];
//       nc                         = rx_phy_postflop_0 [ 164];
//       nc                         = rx_phy_postflop_0 [ 165];
//       nc                         = rx_phy_postflop_0 [ 166];
//       nc                         = rx_phy_postflop_0 [ 167];
//       nc                         = rx_phy_postflop_0 [ 168];
//       nc                         = rx_phy_postflop_0 [ 169];
//       nc                         = rx_phy_postflop_0 [ 170];
//       nc                         = rx_phy_postflop_0 [ 171];
//       nc                         = rx_phy_postflop_0 [ 172];
//       nc                         = rx_phy_postflop_0 [ 173];
//       nc                         = rx_phy_postflop_0 [ 174];
//       nc                         = rx_phy_postflop_0 [ 175];
//       nc                         = rx_phy_postflop_0 [ 176];
//       nc                         = rx_phy_postflop_0 [ 177];
//       nc                         = rx_phy_postflop_0 [ 178];
//       nc                         = rx_phy_postflop_0 [ 179];
//       nc                         = rx_phy_postflop_0 [ 180];
//       nc                         = rx_phy_postflop_0 [ 181];
//       nc                         = rx_phy_postflop_0 [ 182];
//       nc                         = rx_phy_postflop_0 [ 183];
//       nc                         = rx_phy_postflop_0 [ 184];
//       nc                         = rx_phy_postflop_0 [ 185];
//       nc                         = rx_phy_postflop_0 [ 186];
//       nc                         = rx_phy_postflop_0 [ 187];
//       nc                         = rx_phy_postflop_0 [ 188];
//       nc                         = rx_phy_postflop_0 [ 189];
//       nc                         = rx_phy_postflop_0 [ 190];
//       nc                         = rx_phy_postflop_0 [ 191];
//       nc                         = rx_phy_postflop_0 [ 192];
//       nc                         = rx_phy_postflop_0 [ 193];
//       nc                         = rx_phy_postflop_0 [ 194];
//       nc                         = rx_phy_postflop_0 [ 195];
//       nc                         = rx_phy_postflop_0 [ 196];
//       nc                         = rx_phy_postflop_0 [ 197];
//       DBI                        = rx_phy_postflop_0 [ 198];
//       DBI                        = rx_phy_postflop_0 [ 199];
//       nc                         = rx_phy_postflop_0 [ 200];
//       nc                         = rx_phy_postflop_0 [ 201];
//       nc                         = rx_phy_postflop_0 [ 202];
//       nc                         = rx_phy_postflop_0 [ 203];
//       nc                         = rx_phy_postflop_0 [ 204];
//       nc                         = rx_phy_postflop_0 [ 205];
//       nc                         = rx_phy_postflop_0 [ 206];
//       nc                         = rx_phy_postflop_0 [ 207];
//       nc                         = rx_phy_postflop_0 [ 208];
//       nc                         = rx_phy_postflop_0 [ 209];
//       nc                         = rx_phy_postflop_0 [ 210];
//       nc                         = rx_phy_postflop_0 [ 211];
//       nc                         = rx_phy_postflop_0 [ 212];
//       nc                         = rx_phy_postflop_0 [ 213];
//       nc                         = rx_phy_postflop_0 [ 214];
//       nc                         = rx_phy_postflop_0 [ 215];
//       nc                         = rx_phy_postflop_0 [ 216];
//       nc                         = rx_phy_postflop_0 [ 217];
//       nc                         = rx_phy_postflop_0 [ 218];
//       nc                         = rx_phy_postflop_0 [ 219];
//       nc                         = rx_phy_postflop_0 [ 220];
//       nc                         = rx_phy_postflop_0 [ 221];
//       nc                         = rx_phy_postflop_0 [ 222];
//       nc                         = rx_phy_postflop_0 [ 223];
//       nc                         = rx_phy_postflop_0 [ 224];
//       nc                         = rx_phy_postflop_0 [ 225];
//       nc                         = rx_phy_postflop_0 [ 226];
//       nc                         = rx_phy_postflop_0 [ 227];
//       nc                         = rx_phy_postflop_0 [ 228];
//       nc                         = rx_phy_postflop_0 [ 229];
//       nc                         = rx_phy_postflop_0 [ 230];
//       nc                         = rx_phy_postflop_0 [ 231];
//       nc                         = rx_phy_postflop_0 [ 232];
//       nc                         = rx_phy_postflop_0 [ 233];
//       nc                         = rx_phy_postflop_0 [ 234];
//       nc                         = rx_phy_postflop_0 [ 235];
//       nc                         = rx_phy_postflop_0 [ 236];
//       nc                         = rx_phy_postflop_0 [ 237];
//       DBI                        = rx_phy_postflop_0 [ 238];
//       DBI                        = rx_phy_postflop_0 [ 239];
//       MARKER                     = rx_phy_postflop_1 [ 160]
//       STROBE                     = rx_phy_postflop_1 [ 161]
//       nc                         = rx_phy_postflop_1 [ 162];
//       nc                         = rx_phy_postflop_1 [ 163];
//       nc                         = rx_phy_postflop_1 [ 164];
//       nc                         = rx_phy_postflop_1 [ 165];
//       nc                         = rx_phy_postflop_1 [ 166];
//       nc                         = rx_phy_postflop_1 [ 167];
//       nc                         = rx_phy_postflop_1 [ 168];
//       nc                         = rx_phy_postflop_1 [ 169];
//       nc                         = rx_phy_postflop_1 [ 170];
//       nc                         = rx_phy_postflop_1 [ 171];
//       nc                         = rx_phy_postflop_1 [ 172];
//       nc                         = rx_phy_postflop_1 [ 173];
//       nc                         = rx_phy_postflop_1 [ 174];
//       nc                         = rx_phy_postflop_1 [ 175];
//       nc                         = rx_phy_postflop_1 [ 176];
//       nc                         = rx_phy_postflop_1 [ 177];
//       nc                         = rx_phy_postflop_1 [ 178];
//       nc                         = rx_phy_postflop_1 [ 179];
//       nc                         = rx_phy_postflop_1 [ 180];
//       nc                         = rx_phy_postflop_1 [ 181];
//       nc                         = rx_phy_postflop_1 [ 182];
//       nc                         = rx_phy_postflop_1 [ 183];
//       nc                         = rx_phy_postflop_1 [ 184];
//       nc                         = rx_phy_postflop_1 [ 185];
//       nc                         = rx_phy_postflop_1 [ 186];
//       nc                         = rx_phy_postflop_1 [ 187];
//       nc                         = rx_phy_postflop_1 [ 188];
//       nc                         = rx_phy_postflop_1 [ 189];
//       nc                         = rx_phy_postflop_1 [ 190];
//       nc                         = rx_phy_postflop_1 [ 191];
//       nc                         = rx_phy_postflop_1 [ 192];
//       nc                         = rx_phy_postflop_1 [ 193];
//       nc                         = rx_phy_postflop_1 [ 194];
//       nc                         = rx_phy_postflop_1 [ 195];
//       nc                         = rx_phy_postflop_1 [ 196];
//       nc                         = rx_phy_postflop_1 [ 197];
//       DBI                        = rx_phy_postflop_1 [ 198];
//       DBI                        = rx_phy_postflop_1 [ 199];
//       nc                         = rx_phy_postflop_1 [ 200];
//       nc                         = rx_phy_postflop_1 [ 201];
//       nc                         = rx_phy_postflop_1 [ 202];
//       nc                         = rx_phy_postflop_1 [ 203];
//       nc                         = rx_phy_postflop_1 [ 204];
//       nc                         = rx_phy_postflop_1 [ 205];
//       nc                         = rx_phy_postflop_1 [ 206];
//       nc                         = rx_phy_postflop_1 [ 207];
//       nc                         = rx_phy_postflop_1 [ 208];
//       nc                         = rx_phy_postflop_1 [ 209];
//       nc                         = rx_phy_postflop_1 [ 210];
//       nc                         = rx_phy_postflop_1 [ 211];
//       nc                         = rx_phy_postflop_1 [ 212];
//       nc                         = rx_phy_postflop_1 [ 213];
//       nc                         = rx_phy_postflop_1 [ 214];
//       nc                         = rx_phy_postflop_1 [ 215];
//       nc                         = rx_phy_postflop_1 [ 216];
//       nc                         = rx_phy_postflop_1 [ 217];
//       nc                         = rx_phy_postflop_1 [ 218];
//       nc                         = rx_phy_postflop_1 [ 219];
//       nc                         = rx_phy_postflop_1 [ 220];
//       nc                         = rx_phy_postflop_1 [ 221];
//       nc                         = rx_phy_postflop_1 [ 222];
//       nc                         = rx_phy_postflop_1 [ 223];
//       nc                         = rx_phy_postflop_1 [ 224];
//       nc                         = rx_phy_postflop_1 [ 225];
//       nc                         = rx_phy_postflop_1 [ 226];
//       nc                         = rx_phy_postflop_1 [ 227];
//       nc                         = rx_phy_postflop_1 [ 228];
//       nc                         = rx_phy_postflop_1 [ 229];
//       nc                         = rx_phy_postflop_1 [ 230];
//       nc                         = rx_phy_postflop_1 [ 231];
//       nc                         = rx_phy_postflop_1 [ 232];
//       nc                         = rx_phy_postflop_1 [ 233];
//       nc                         = rx_phy_postflop_1 [ 234];
//       nc                         = rx_phy_postflop_1 [ 235];
//       nc                         = rx_phy_postflop_1 [ 236];
//       nc                         = rx_phy_postflop_1 [ 237];
//       DBI                        = rx_phy_postflop_1 [ 238];
//       DBI                        = rx_phy_postflop_1 [ 239];
//       MARKER                     = rx_phy_postflop_0 [ 240]
//       STROBE                     = rx_phy_postflop_0 [ 241]
  assign rx_st_credit_r3            = rx_phy_postflop_0 [ 242];
//       nc                         = rx_phy_postflop_0 [ 243];
//       nc                         = rx_phy_postflop_0 [ 244];
//       nc                         = rx_phy_postflop_0 [ 245];
//       nc                         = rx_phy_postflop_0 [ 246];
//       nc                         = rx_phy_postflop_0 [ 247];
//       nc                         = rx_phy_postflop_0 [ 248];
//       nc                         = rx_phy_postflop_0 [ 249];
//       nc                         = rx_phy_postflop_0 [ 250];
//       nc                         = rx_phy_postflop_0 [ 251];
//       nc                         = rx_phy_postflop_0 [ 252];
//       nc                         = rx_phy_postflop_0 [ 253];
//       nc                         = rx_phy_postflop_0 [ 254];
//       nc                         = rx_phy_postflop_0 [ 255];
//       nc                         = rx_phy_postflop_0 [ 256];
//       nc                         = rx_phy_postflop_0 [ 257];
//       nc                         = rx_phy_postflop_0 [ 258];
//       nc                         = rx_phy_postflop_0 [ 259];
//       nc                         = rx_phy_postflop_0 [ 260];
//       nc                         = rx_phy_postflop_0 [ 261];
//       nc                         = rx_phy_postflop_0 [ 262];
//       nc                         = rx_phy_postflop_0 [ 263];
//       nc                         = rx_phy_postflop_0 [ 264];
//       nc                         = rx_phy_postflop_0 [ 265];
//       nc                         = rx_phy_postflop_0 [ 266];
//       nc                         = rx_phy_postflop_0 [ 267];
//       nc                         = rx_phy_postflop_0 [ 268];
//       nc                         = rx_phy_postflop_0 [ 269];
//       nc                         = rx_phy_postflop_0 [ 270];
//       nc                         = rx_phy_postflop_0 [ 271];
//       nc                         = rx_phy_postflop_0 [ 272];
//       nc                         = rx_phy_postflop_0 [ 273];
//       nc                         = rx_phy_postflop_0 [ 274];
//       nc                         = rx_phy_postflop_0 [ 275];
//       nc                         = rx_phy_postflop_0 [ 276];
//       nc                         = rx_phy_postflop_0 [ 277];
//       DBI                        = rx_phy_postflop_0 [ 278];
//       DBI                        = rx_phy_postflop_0 [ 279];
//       nc                         = rx_phy_postflop_0 [ 280];
//       nc                         = rx_phy_postflop_0 [ 281];
//       nc                         = rx_phy_postflop_0 [ 282];
//       nc                         = rx_phy_postflop_0 [ 283];
//       nc                         = rx_phy_postflop_0 [ 284];
//       nc                         = rx_phy_postflop_0 [ 285];
//       nc                         = rx_phy_postflop_0 [ 286];
//       nc                         = rx_phy_postflop_0 [ 287];
//       nc                         = rx_phy_postflop_0 [ 288];
//       nc                         = rx_phy_postflop_0 [ 289];
//       nc                         = rx_phy_postflop_0 [ 290];
//       nc                         = rx_phy_postflop_0 [ 291];
//       nc                         = rx_phy_postflop_0 [ 292];
//       nc                         = rx_phy_postflop_0 [ 293];
//       nc                         = rx_phy_postflop_0 [ 294];
//       nc                         = rx_phy_postflop_0 [ 295];
//       nc                         = rx_phy_postflop_0 [ 296];
//       nc                         = rx_phy_postflop_0 [ 297];
//       nc                         = rx_phy_postflop_0 [ 298];
//       nc                         = rx_phy_postflop_0 [ 299];
//       nc                         = rx_phy_postflop_0 [ 300];
//       nc                         = rx_phy_postflop_0 [ 301];
//       nc                         = rx_phy_postflop_0 [ 302];
//       nc                         = rx_phy_postflop_0 [ 303];
//       nc                         = rx_phy_postflop_0 [ 304];
//       nc                         = rx_phy_postflop_0 [ 305];
//       nc                         = rx_phy_postflop_0 [ 306];
//       nc                         = rx_phy_postflop_0 [ 307];
//       nc                         = rx_phy_postflop_0 [ 308];
//       nc                         = rx_phy_postflop_0 [ 309];
//       nc                         = rx_phy_postflop_0 [ 310];
//       nc                         = rx_phy_postflop_0 [ 311];
//       nc                         = rx_phy_postflop_0 [ 312];
//       nc                         = rx_phy_postflop_0 [ 313];
//       nc                         = rx_phy_postflop_0 [ 314];
//       nc                         = rx_phy_postflop_0 [ 315];
//       nc                         = rx_phy_postflop_0 [ 316];
//       nc                         = rx_phy_postflop_0 [ 317];
//       DBI                        = rx_phy_postflop_0 [ 318];
//       DBI                        = rx_phy_postflop_0 [ 319];
//       MARKER                     = rx_phy_postflop_1 [ 240]
//       STROBE                     = rx_phy_postflop_1 [ 241]
//       nc                         = rx_phy_postflop_1 [ 242];
//       nc                         = rx_phy_postflop_1 [ 243];
//       nc                         = rx_phy_postflop_1 [ 244];
//       nc                         = rx_phy_postflop_1 [ 245];
//       nc                         = rx_phy_postflop_1 [ 246];
//       nc                         = rx_phy_postflop_1 [ 247];
//       nc                         = rx_phy_postflop_1 [ 248];
//       nc                         = rx_phy_postflop_1 [ 249];
//       nc                         = rx_phy_postflop_1 [ 250];
//       nc                         = rx_phy_postflop_1 [ 251];
//       nc                         = rx_phy_postflop_1 [ 252];
//       nc                         = rx_phy_postflop_1 [ 253];
//       nc                         = rx_phy_postflop_1 [ 254];
//       nc                         = rx_phy_postflop_1 [ 255];
//       nc                         = rx_phy_postflop_1 [ 256];
//       nc                         = rx_phy_postflop_1 [ 257];
//       nc                         = rx_phy_postflop_1 [ 258];
//       nc                         = rx_phy_postflop_1 [ 259];
//       nc                         = rx_phy_postflop_1 [ 260];
//       nc                         = rx_phy_postflop_1 [ 261];
//       nc                         = rx_phy_postflop_1 [ 262];
//       nc                         = rx_phy_postflop_1 [ 263];
//       nc                         = rx_phy_postflop_1 [ 264];
//       nc                         = rx_phy_postflop_1 [ 265];
//       nc                         = rx_phy_postflop_1 [ 266];
//       nc                         = rx_phy_postflop_1 [ 267];
//       nc                         = rx_phy_postflop_1 [ 268];
//       nc                         = rx_phy_postflop_1 [ 269];
//       nc                         = rx_phy_postflop_1 [ 270];
//       nc                         = rx_phy_postflop_1 [ 271];
//       nc                         = rx_phy_postflop_1 [ 272];
//       nc                         = rx_phy_postflop_1 [ 273];
//       nc                         = rx_phy_postflop_1 [ 274];
//       nc                         = rx_phy_postflop_1 [ 275];
//       nc                         = rx_phy_postflop_1 [ 276];
//       nc                         = rx_phy_postflop_1 [ 277];
//       DBI                        = rx_phy_postflop_1 [ 278];
//       DBI                        = rx_phy_postflop_1 [ 279];
//       nc                         = rx_phy_postflop_1 [ 280];
//       nc                         = rx_phy_postflop_1 [ 281];
//       nc                         = rx_phy_postflop_1 [ 282];
//       nc                         = rx_phy_postflop_1 [ 283];
//       nc                         = rx_phy_postflop_1 [ 284];
//       nc                         = rx_phy_postflop_1 [ 285];
//       nc                         = rx_phy_postflop_1 [ 286];
//       nc                         = rx_phy_postflop_1 [ 287];
//       nc                         = rx_phy_postflop_1 [ 288];
//       nc                         = rx_phy_postflop_1 [ 289];
//       nc                         = rx_phy_postflop_1 [ 290];
//       nc                         = rx_phy_postflop_1 [ 291];
//       nc                         = rx_phy_postflop_1 [ 292];
//       nc                         = rx_phy_postflop_1 [ 293];
//       nc                         = rx_phy_postflop_1 [ 294];
//       nc                         = rx_phy_postflop_1 [ 295];
//       nc                         = rx_phy_postflop_1 [ 296];
//       nc                         = rx_phy_postflop_1 [ 297];
//       nc                         = rx_phy_postflop_1 [ 298];
//       nc                         = rx_phy_postflop_1 [ 299];
//       nc                         = rx_phy_postflop_1 [ 300];
//       nc                         = rx_phy_postflop_1 [ 301];
//       nc                         = rx_phy_postflop_1 [ 302];
//       nc                         = rx_phy_postflop_1 [ 303];
//       nc                         = rx_phy_postflop_1 [ 304];
//       nc                         = rx_phy_postflop_1 [ 305];
//       nc                         = rx_phy_postflop_1 [ 306];
//       nc                         = rx_phy_postflop_1 [ 307];
//       nc                         = rx_phy_postflop_1 [ 308];
//       nc                         = rx_phy_postflop_1 [ 309];
//       nc                         = rx_phy_postflop_1 [ 310];
//       nc                         = rx_phy_postflop_1 [ 311];
//       nc                         = rx_phy_postflop_1 [ 312];
//       nc                         = rx_phy_postflop_1 [ 313];
//       nc                         = rx_phy_postflop_1 [ 314];
//       nc                         = rx_phy_postflop_1 [ 315];
//       nc                         = rx_phy_postflop_1 [ 316];
//       nc                         = rx_phy_postflop_1 [ 317];
//       DBI                        = rx_phy_postflop_1 [ 318];
//       DBI                        = rx_phy_postflop_1 [ 319];

// RX Section
//////////////////////////////////////////////////////////////////


endmodule
